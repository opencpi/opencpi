-- This package enables VHDL code to instantiate all entities and modules in this library
library ieee; use IEEE.std_logic_1164.all; use ieee.numeric_std.all;
library ocpi; use ocpi.types.all;
library platform; use platform.platform_pkg.all;
library axi; use axi.axi_pkg.all;
package zynq_ultra_pkg is

-- Signals from the PS for use by the PL
type ps2pl_t is record
  FCLK         : std_logic_vector(3 downto 0);
  FCLKRESET_N  : std_logic;
end record ps2pl_t;
-- Signals from the PL for use by the PS
type pl2ps_t is record
  DEBUG        : std_logic_vector(31 downto 0); --     FTMT_F2P_DEBUG
end record pl2ps_t;


component zynq_ultra_ps_e_v3_2_1 is
  generic (
    C_MAXIGP0_DATA_WIDTH : integer := 32;
    C_MAXIGP1_DATA_WIDTH : integer := 32;
    C_MAXIGP2_DATA_WIDTH : integer := 128;

    C_SAXIGP0_DATA_WIDTH : integer := 128;
    C_SAXIGP1_DATA_WIDTH : integer := 128;
    C_SAXIGP2_DATA_WIDTH : integer := 64;
    C_SAXIGP3_DATA_WIDTH : integer := 64;
    C_SAXIGP4_DATA_WIDTH : integer := 64;
    C_SAXIGP5_DATA_WIDTH : integer := 64;
    C_SAXIGP6_DATA_WIDTH : integer := 128;
    C_SD0_INTERNAL_BUS_WIDTH : integer := 8;
    C_SD1_INTERNAL_BUS_WIDTH : integer := 8;
    C_PL_CLK0_BUF : string := "TRUE";
    C_PL_CLK1_BUF : string := "TRUE";
    C_PL_CLK2_BUF : string := "TRUE";
    C_PL_CLK3_BUF : string := "TRUE";

    C_NUM_F2P_0_INTR_INPUTS : integer := 0;
    C_NUM_F2P_1_INTR_INPUTS : integer := 0;

    C_NUM_FABRIC_RESETS : integer := 1;
    C_EMIO_GPIO_WIDTH : integer := 64; -- was 96

--    C_TRISTATE_INVERTED : integer := 1;

    C_USE_DIFF_RW_CLK_GP0 : integer := 0;
    C_USE_DIFF_RW_CLK_GP1 : integer := 0;
    C_USE_DIFF_RW_CLK_GP2 : integer := 0;
    C_USE_DIFF_RW_CLK_GP3 : integer := 0;
    C_USE_DIFF_RW_CLK_GP4 : integer := 0;
    C_USE_DIFF_RW_CLK_GP5 : integer := 0;
    C_USE_DIFF_RW_CLK_GP6 : integer := 0;

    C_TRACE_PIPELINE_WIDTH : integer := 8;
    C_EN_EMIO_TRACE : integer := 0;
    C_EN_FIFO_ENET0 : integer := 0;
    C_EN_FIFO_ENET1 : integer := 0;
    C_EN_FIFO_ENET2 : integer := 0;
    C_EN_FIFO_ENET3 : integer := 0;
    C_TRACE_DATA_WIDTH : integer := 32;

    C_USE_DEBUG_TEST : integer := 0;
    C_DP_USE_AUDIO : integer := 0;
    C_DP_USE_VIDEO : integer := 0
);
  port (
-- maxigp0
    maxihpm0_fpd_aclk : in std_logic;
    dp_video_ref_clk : out std_logic;
    dp_audio_ref_clk : out std_logic;
    maxigp0_awid : out std_logic_vector(15 downto 0);
    maxigp0_awaddr : out std_logic_vector(39 downto 0);
    maxigp0_awlen : out std_logic_vector(7 downto 0);
    maxigp0_awsize : out std_logic_vector(2 downto 0);
    maxigp0_awburst : out std_logic_vector(1 downto 0);
    maxigp0_awlock : out std_logic;
    maxigp0_awcache : out std_logic_vector(3 downto 0);
    maxigp0_awprot : out std_logic_vector(2 downto 0);
    maxigp0_awvalid : out std_logic;
    maxigp0_awuser : out std_logic_vector(15 downto 0);
    maxigp0_awready : in std_logic;
    maxigp0_wdata : out std_logic_vector(C_MAXIGP0_DATA_WIDTH-1  downto 0);
    maxigp0_wstrb : out std_logic_vector((C_MAXIGP0_DATA_WIDTH/8)-1  downto 0);
    maxigp0_wlast : out std_logic;
    maxigp0_wvalid : out std_logic;
    maxigp0_wready : in std_logic;
    maxigp0_bid : in std_logic_vector(15 downto 0);
    maxigp0_bresp : in std_logic_vector(1 downto 0);
    maxigp0_bvalid : in std_logic;
    maxigp0_bready : out std_logic;
    maxigp0_arid : out std_logic_vector(15 downto 0);
    maxigp0_araddr : out std_logic_vector(39 downto 0);
    maxigp0_arlen : out std_logic_vector(7 downto 0);
    maxigp0_arsize : out std_logic_vector(2 downto 0);
    maxigp0_arburst : out std_logic_vector(1 downto 0);
    maxigp0_arlock : out std_logic;
    maxigp0_arcache : out std_logic_vector(3 downto 0);
    maxigp0_arprot : out std_logic_vector(2 downto 0);
    maxigp0_arvalid : out std_logic;
    maxigp0_aruser : out std_logic_vector(15 downto 0);
    maxigp0_arready : in std_logic;
    maxigp0_rid : in std_logic_vector(15 downto 0);
    maxigp0_rdata : in std_logic_vector(C_MAXIGP0_DATA_WIDTH-1  downto 0);
    maxigp0_rresp : in std_logic_vector(1 downto 0);
    maxigp0_rlast : in std_logic;
    maxigp0_rvalid : in std_logic;
    maxigp0_rready : out std_logic;
    maxigp0_awqos : out std_logic_vector(3 downto 0);
    maxigp0_arqos : out std_logic_vector(3 downto 0);

-- maxigp1
    maxihpm1_fpd_aclk : in std_logic;
    maxigp1_awid : out std_logic_vector(15 downto 0);
    maxigp1_awaddr : out std_logic_vector(39 downto 0);
    maxigp1_awlen : out std_logic_vector(7 downto 0);
    maxigp1_awsize : out std_logic_vector(2 downto 0);
    maxigp1_awburst : out std_logic_vector(1 downto 0);
    maxigp1_awlock : out std_logic;
    maxigp1_awcache : out std_logic_vector(3 downto 0);
    maxigp1_awprot : out std_logic_vector(2 downto 0);
    maxigp1_awvalid : out std_logic;
    maxigp1_awuser : out std_logic_vector(15 downto 0);
    maxigp1_awready : in std_logic;
    maxigp1_wdata : out std_logic_vector(C_MAXIGP1_DATA_WIDTH-1  downto 0);
    maxigp1_wstrb : out std_logic_vector((C_MAXIGP1_DATA_WIDTH/8)-1  downto 0);
    maxigp1_wlast : out std_logic;
    maxigp1_wvalid : out std_logic;
    maxigp1_wready : in std_logic;
    maxigp1_bid : in std_logic_vector(15 downto 0);
    maxigp1_bresp : in std_logic_vector(1 downto 0);
    maxigp1_bvalid : in std_logic;
    maxigp1_bready : out std_logic;
    maxigp1_arid : out std_logic_vector(15 downto 0);
    maxigp1_araddr : out std_logic_vector(39 downto 0);
    maxigp1_arlen : out std_logic_vector(7 downto 0);
    maxigp1_arsize : out std_logic_vector(2 downto 0);
    maxigp1_arburst : out std_logic_vector(1 downto 0);
    maxigp1_arlock : out std_logic;
    maxigp1_arcache : out std_logic_vector(3 downto 0);
    maxigp1_arprot : out std_logic_vector(2 downto 0);
    maxigp1_arvalid : out std_logic;
    maxigp1_aruser : out std_logic_vector(15 downto 0);
    maxigp1_arready : in std_logic;
    maxigp1_rid : in std_logic_vector(15 downto 0);
    maxigp1_rdata : in std_logic_vector(C_MAXIGP1_DATA_WIDTH-1  downto 0);
    maxigp1_rresp : in std_logic_vector(1 downto 0);
    maxigp1_rlast : in std_logic;
    maxigp1_rvalid : in std_logic;
    maxigp1_rready : out std_logic;
    maxigp1_awqos : out std_logic_vector(3 downto 0);
    maxigp1_arqos : out std_logic_vector(3 downto 0);
-- maxigp2
    maxihpm0_lpd_aclk : in std_logic;
    maxigp2_awid : out std_logic_vector(15 downto 0);
    maxigp2_awaddr : out std_logic_vector(39 downto 0);
    maxigp2_awlen : out std_logic_vector(7 downto 0);
    maxigp2_awsize : out std_logic_vector(2 downto 0);
    maxigp2_awburst : out std_logic_vector(1 downto 0);
    maxigp2_awlock : out std_logic;
    maxigp2_awcache : out std_logic_vector(3 downto 0);
    maxigp2_awprot : out std_logic_vector(2 downto 0);
    maxigp2_awvalid : out std_logic;
    maxigp2_awuser : out std_logic_vector(15 downto 0);
    maxigp2_awready : in std_logic;
    maxigp2_wdata : out std_logic_vector(C_MAXIGP2_DATA_WIDTH-1  downto 0);
    maxigp2_wstrb : out std_logic_vector((C_MAXIGP2_DATA_WIDTH/8)-1  downto 0);
    maxigp2_wlast : out std_logic;
    maxigp2_wvalid : out std_logic;
    maxigp2_wready : in std_logic;
    maxigp2_bid : in std_logic_vector(15 downto 0);
    maxigp2_bresp : in std_logic_vector(1 downto 0);
    maxigp2_bvalid : in std_logic;
    maxigp2_bready : out std_logic;
    maxigp2_arid : out std_logic_vector(15 downto 0);
    maxigp2_araddr : out std_logic_vector(39 downto 0);
    maxigp2_arlen : out std_logic_vector(7 downto 0);
    maxigp2_arsize : out std_logic_vector(2 downto 0);
    maxigp2_arburst : out std_logic_vector(1 downto 0);
    maxigp2_arlock : out std_logic;
    maxigp2_arcache : out std_logic_vector(3 downto 0);
    maxigp2_arprot : out std_logic_vector(2 downto 0);
    maxigp2_arvalid : out std_logic;
    maxigp2_aruser : out std_logic_vector(15 downto 0);
    maxigp2_arready : in std_logic;
    maxigp2_rid : in std_logic_vector(15 downto 0);
    maxigp2_rdata : in std_logic_vector(C_MAXIGP2_DATA_WIDTH-1  downto 0);
    maxigp2_rresp : in std_logic_vector(1 downto 0);
    maxigp2_rlast : in std_logic;
    maxigp2_rvalid : in std_logic;
    maxigp2_rready : out std_logic;
    maxigp2_awqos : out std_logic_vector(3 downto 0);
    maxigp2_arqos : out std_logic_vector(3 downto 0);
-- saxigp0
    saxihpc0_fpd_aclk : in std_logic;
    saxihpc0_fpd_rclk : in std_logic;
    saxihpc0_fpd_wclk : in std_logic;
    saxigp0_aruser : in std_logic;
    saxigp0_awuser : in std_logic;
    saxigp0_awid : in std_logic_vector(5 downto 0);
    saxigp0_awaddr : in std_logic_vector(48 downto 0);
    saxigp0_awlen : in std_logic_vector(7 downto 0);
    saxigp0_awsize : in std_logic_vector(2 downto 0);
    saxigp0_awburst : in std_logic_vector(1 downto 0);
    saxigp0_awlock : in std_logic;
    saxigp0_awcache : in std_logic_vector(3 downto 0);
    saxigp0_awprot : in std_logic_vector(2 downto 0);
    saxigp0_awvalid : in std_logic;
    saxigp0_awready : out std_logic;
    saxigp0_wdata : in std_logic_vector(C_SAXIGP0_DATA_WIDTH-1 downto 0);
    saxigp0_wstrb : in std_logic_vector((C_SAXIGP0_DATA_WIDTH/8) -1  downto 0);
    saxigp0_wlast : in std_logic;
    saxigp0_wvalid : in std_logic;
    saxigp0_wready : out std_logic;
    saxigp0_bid : out std_logic_vector(5 downto 0);
    saxigp0_bresp : out std_logic_vector(1 downto 0);
    saxigp0_bvalid : out std_logic;
    saxigp0_bready : in std_logic;
    saxigp0_arid : in std_logic_vector(5 downto 0);
    saxigp0_araddr : in std_logic_vector(48 downto 0);
    saxigp0_arlen : in std_logic_vector(7 downto 0);
    saxigp0_arsize : in std_logic_vector(2 downto 0);
    saxigp0_arburst : in std_logic_vector(1 downto 0);
    saxigp0_arlock : in std_logic;
    saxigp0_arcache : in std_logic_vector(3 downto 0);
    saxigp0_arprot : in std_logic_vector(2 downto 0);
    saxigp0_arvalid : in std_logic;
    saxigp0_arready : out std_logic;
    saxigp0_rid : out std_logic_vector(5 downto 0);
    saxigp0_rdata : out std_logic_vector(C_SAXIGP0_DATA_WIDTH-1 downto 0);
    saxigp0_rresp : out std_logic_vector(1 downto 0);
    saxigp0_rlast : out std_logic;
    saxigp0_rvalid : out std_logic;
    saxigp0_rready : in std_logic;
    saxigp0_awqos : in std_logic_vector(3 downto 0);
    saxigp0_arqos : in std_logic_vector(3 downto 0);
    saxigp0_rcount : out std_logic_vector(7 downto 0);
    saxigp0_wcount : out std_logic_vector(7 downto 0);
    saxigp0_racount : out std_logic_vector(3 downto 0);
    saxigp0_wacount : out std_logic_vector(3 downto 0);
-- saxigp1
    saxihpc1_fpd_aclk : in std_logic;
    saxihpc1_fpd_rclk : in std_logic;
    saxihpc1_fpd_wclk : in std_logic;
    saxigp1_aruser : in std_logic;
    saxigp1_awuser : in std_logic;
    saxigp1_awid : in std_logic_vector(5 downto 0);
    saxigp1_awaddr : in std_logic_vector(48 downto 0);
    saxigp1_awlen : in std_logic_vector(7 downto 0);
    saxigp1_awsize : in std_logic_vector(2 downto 0);
    saxigp1_awburst : in std_logic_vector(1 downto 0);
    saxigp1_awlock : in std_logic;
    saxigp1_awcache : in std_logic_vector(3 downto 0);
    saxigp1_awprot : in std_logic_vector(2 downto 0);
    saxigp1_awvalid : in std_logic;
    saxigp1_awready : out std_logic;
    saxigp1_wdata : in std_logic_vector(C_SAXIGP1_DATA_WIDTH-1 downto 0);
    saxigp1_wstrb : in std_logic_vector((C_SAXIGP1_DATA_WIDTH/8) -1  downto 0);
    saxigp1_wlast : in std_logic;
    saxigp1_wvalid : in std_logic;
    saxigp1_wready : out std_logic;
    saxigp1_bid : out std_logic_vector(5 downto 0);
    saxigp1_bresp : out std_logic_vector(1 downto 0);
    saxigp1_bvalid : out std_logic;
    saxigp1_bready : in std_logic;
    saxigp1_arid : in std_logic_vector(5 downto 0);
    saxigp1_araddr : in std_logic_vector(48 downto 0);
    saxigp1_arlen : in std_logic_vector(7 downto 0);
    saxigp1_arsize : in std_logic_vector(2 downto 0);
    saxigp1_arburst : in std_logic_vector(1 downto 0);
    saxigp1_arlock : in std_logic;
    saxigp1_arcache : in std_logic_vector(3 downto 0);
    saxigp1_arprot : in std_logic_vector(2 downto 0);
    saxigp1_arvalid : in std_logic;
    saxigp1_arready : out std_logic;
    saxigp1_rid : out std_logic_vector(5 downto 0);
    saxigp1_rdata : out std_logic_vector(C_SAXIGP1_DATA_WIDTH-1 downto 0);
    saxigp1_rresp : out std_logic_vector(1 downto 0);
    saxigp1_rlast : out std_logic;
    saxigp1_rvalid : out std_logic;
    saxigp1_rready : in std_logic;
    saxigp1_awqos : in std_logic_vector(3 downto 0);
    saxigp1_arqos : in std_logic_vector(3 downto 0);
    saxigp1_rcount : out std_logic_vector(7 downto 0);
    saxigp1_wcount : out std_logic_vector(7 downto 0);
    saxigp1_racount : out std_logic_vector(3 downto 0);
    saxigp1_wacount : out std_logic_vector(3 downto 0);
-- saxigp2
    saxihp0_fpd_aclk : in std_logic;
    saxihp0_fpd_rclk : in std_logic;
    saxihp0_fpd_wclk : in std_logic;
    saxigp2_aruser : in std_logic;
    saxigp2_awuser : in std_logic;
    saxigp2_awid : in std_logic_vector(5 downto 0);
    saxigp2_awaddr : in std_logic_vector(48 downto 0);
    saxigp2_awlen : in std_logic_vector(7 downto 0);
    saxigp2_awsize : in std_logic_vector(2 downto 0);
    saxigp2_awburst : in std_logic_vector(1 downto 0);
    saxigp2_awlock : in std_logic;
    saxigp2_awcache : in std_logic_vector(3 downto 0);
    saxigp2_awprot : in std_logic_vector(2 downto 0);
    saxigp2_awvalid : in std_logic;
    saxigp2_awready : out std_logic;
    saxigp2_wdata : in std_logic_vector(C_SAXIGP2_DATA_WIDTH-1 downto 0);
    saxigp2_wstrb : in std_logic_vector((C_SAXIGP2_DATA_WIDTH/8) -1  downto 0);
    saxigp2_wlast : in std_logic;
    saxigp2_wvalid : in std_logic;
    saxigp2_wready : out std_logic;
    saxigp2_bid : out std_logic_vector(5 downto 0);
    saxigp2_bresp : out std_logic_vector(1 downto 0);
    saxigp2_bvalid : out std_logic;
    saxigp2_bready : in std_logic;
    saxigp2_arid : in std_logic_vector(5 downto 0);
    saxigp2_araddr : in std_logic_vector(48 downto 0);
    saxigp2_arlen : in std_logic_vector(7 downto 0);
    saxigp2_arsize : in std_logic_vector(2 downto 0);
    saxigp2_arburst : in std_logic_vector(1 downto 0);
    saxigp2_arlock : in std_logic;
    saxigp2_arcache : in std_logic_vector(3 downto 0);
    saxigp2_arprot : in std_logic_vector(2 downto 0);
    saxigp2_arvalid : in std_logic;
    saxigp2_arready : out std_logic;
    saxigp2_rid : out std_logic_vector(5 downto 0);
    saxigp2_rdata : out std_logic_vector(C_SAXIGP2_DATA_WIDTH-1 downto 0);
    saxigp2_rresp : out std_logic_vector(1 downto 0);
    saxigp2_rlast : out std_logic;
    saxigp2_rvalid : out std_logic;
    saxigp2_rready : in std_logic;
    saxigp2_awqos : in std_logic_vector(3 downto 0);
    saxigp2_arqos : in std_logic_vector(3 downto 0);
    saxigp2_rcount : out std_logic_vector(7 downto 0);
    saxigp2_wcount : out std_logic_vector(7 downto 0);
    saxigp2_racount : out std_logic_vector(3 downto 0);
    saxigp2_wacount : out std_logic_vector(3 downto 0);
-- saxigp3
    saxihp1_fpd_aclk : in std_logic;
    saxihp1_fpd_rclk : in std_logic;
    saxihp1_fpd_wclk : in std_logic;
    saxigp3_aruser : in std_logic;
    saxigp3_awuser : in std_logic;
    saxigp3_awid : in std_logic_vector(5 downto 0);
    saxigp3_awaddr : in std_logic_vector(48 downto 0);
    saxigp3_awlen : in std_logic_vector(7 downto 0);
    saxigp3_awsize : in std_logic_vector(2 downto 0);
    saxigp3_awburst : in std_logic_vector(1 downto 0);
    saxigp3_awlock : in std_logic;
    saxigp3_awcache : in std_logic_vector(3 downto 0);
    saxigp3_awprot : in std_logic_vector(2 downto 0);
    saxigp3_awvalid : in std_logic;
    saxigp3_awready : out std_logic;
    saxigp3_wdata : in std_logic_vector(C_SAXIGP3_DATA_WIDTH-1 downto 0);
    saxigp3_wstrb : in std_logic_vector((C_SAXIGP3_DATA_WIDTH/8) -1  downto 0);
    saxigp3_wlast : in std_logic;
    saxigp3_wvalid : in std_logic;
    saxigp3_wready : out std_logic;
    saxigp3_bid : out std_logic_vector(5 downto 0);
    saxigp3_bresp : out std_logic_vector(1 downto 0);
    saxigp3_bvalid : out std_logic;
    saxigp3_bready : in std_logic;
    saxigp3_arid : in std_logic_vector(5 downto 0);
    saxigp3_araddr : in std_logic_vector(48 downto 0);
    saxigp3_arlen : in std_logic_vector(7 downto 0);
    saxigp3_arsize : in std_logic_vector(2 downto 0);
    saxigp3_arburst : in std_logic_vector(1 downto 0);
    saxigp3_arlock : in std_logic;
    saxigp3_arcache : in std_logic_vector(3 downto 0);
    saxigp3_arprot : in std_logic_vector(2 downto 0);
    saxigp3_arvalid : in std_logic;
    saxigp3_arready : out std_logic;
    saxigp3_rid : out std_logic_vector(5 downto 0);
    saxigp3_rdata : out std_logic_vector(C_SAXIGP3_DATA_WIDTH-1 downto 0);
    saxigp3_rresp : out std_logic_vector(1 downto 0);
    saxigp3_rlast : out std_logic;
    saxigp3_rvalid : out std_logic;
    saxigp3_rready : in std_logic;
    saxigp3_awqos : in std_logic_vector(3 downto 0);
    saxigp3_arqos : in std_logic_vector(3 downto 0);
    saxigp3_rcount : out std_logic_vector(7 downto 0);
    saxigp3_wcount : out std_logic_vector(7 downto 0);
    saxigp3_racount : out std_logic_vector(3 downto 0);
    saxigp3_wacount : out std_logic_vector(3 downto 0);
-- saxigp4
    saxihp2_fpd_aclk : in std_logic;
    saxihp2_fpd_rclk : in std_logic;
    saxihp2_fpd_wclk : in std_logic;
    saxigp4_aruser : in std_logic;
    saxigp4_awuser : in std_logic;
    saxigp4_awid : in std_logic_vector(5 downto 0);
    saxigp4_awaddr : in std_logic_vector(48 downto 0);
    saxigp4_awlen : in std_logic_vector(7 downto 0);
    saxigp4_awsize : in std_logic_vector(2 downto 0);
    saxigp4_awburst : in std_logic_vector(1 downto 0);
    saxigp4_awlock : in std_logic;
    saxigp4_awcache : in std_logic_vector(3 downto 0);
    saxigp4_awprot : in std_logic_vector(2 downto 0);
    saxigp4_awvalid : in std_logic;
    saxigp4_awready : out std_logic;
    saxigp4_wdata : in std_logic_vector(C_SAXIGP4_DATA_WIDTH-1 downto 0);
    saxigp4_wstrb : in std_logic_vector((C_SAXIGP4_DATA_WIDTH/8) -1  downto 0);
    saxigp4_wlast : in std_logic;
    saxigp4_wvalid : in std_logic;
    saxigp4_wready : out std_logic;
    saxigp4_bid : out std_logic_vector(5 downto 0);
    saxigp4_bresp : out std_logic_vector(1 downto 0);
    saxigp4_bvalid : out std_logic;
    saxigp4_bready : in std_logic;
    saxigp4_arid : in std_logic_vector(5 downto 0);
    saxigp4_araddr : in std_logic_vector(48 downto 0);
    saxigp4_arlen : in std_logic_vector(7 downto 0);
    saxigp4_arsize : in std_logic_vector(2 downto 0);
    saxigp4_arburst : in std_logic_vector(1 downto 0);
    saxigp4_arlock : in std_logic;
    saxigp4_arcache : in std_logic_vector(3 downto 0);
    saxigp4_arprot : in std_logic_vector(2 downto 0);
    saxigp4_arvalid : in std_logic;
    saxigp4_arready : out std_logic;
    saxigp4_rid : out std_logic_vector(5 downto 0);
    saxigp4_rdata : out std_logic_vector(C_SAXIGP4_DATA_WIDTH-1 downto 0);
    saxigp4_rresp : out std_logic_vector(1 downto 0);
    saxigp4_rlast : out std_logic;
    saxigp4_rvalid : out std_logic;
    saxigp4_rready : in std_logic;
    saxigp4_awqos : in std_logic_vector(3 downto 0);
    saxigp4_arqos : in std_logic_vector(3 downto 0);
    saxigp4_rcount : out std_logic_vector(7 downto 0);
    saxigp4_wcount : out std_logic_vector(7 downto 0);
    saxigp4_racount : out std_logic_vector(3 downto 0);
    saxigp4_wacount : out std_logic_vector(3 downto 0);
-- saxigp5
    saxihp3_fpd_aclk : in std_logic;
    saxihp3_fpd_rclk : in std_logic;
    saxihp3_fpd_wclk : in std_logic;
    saxigp5_aruser : in std_logic;
    saxigp5_awuser : in std_logic;
    saxigp5_awid : in std_logic_vector(5 downto 0);
    saxigp5_awaddr : in std_logic_vector(48 downto 0);
    saxigp5_awlen : in std_logic_vector(7 downto 0);
    saxigp5_awsize : in std_logic_vector(2 downto 0);
    saxigp5_awburst : in std_logic_vector(1 downto 0);
    saxigp5_awlock : in std_logic;
    saxigp5_awcache : in std_logic_vector(3 downto 0);
    saxigp5_awprot : in std_logic_vector(2 downto 0);
    saxigp5_awvalid : in std_logic;
    saxigp5_awready : out std_logic;
    saxigp5_wdata : in std_logic_vector(C_SAXIGP5_DATA_WIDTH-1 downto 0);
    saxigp5_wstrb : in std_logic_vector((C_SAXIGP5_DATA_WIDTH/8) -1  downto 0);
    saxigp5_wlast : in std_logic;
    saxigp5_wvalid : in std_logic;
    saxigp5_wready : out std_logic;
    saxigp5_bid : out std_logic_vector(5 downto 0);
    saxigp5_bresp : out std_logic_vector(1 downto 0);
    saxigp5_bvalid : out std_logic;
    saxigp5_bready : in std_logic;
    saxigp5_arid : in std_logic_vector(5 downto 0);
    saxigp5_araddr : in std_logic_vector(48 downto 0);
    saxigp5_arlen : in std_logic_vector(7 downto 0);
    saxigp5_arsize : in std_logic_vector(2 downto 0);
    saxigp5_arburst : in std_logic_vector(1 downto 0);
    saxigp5_arlock : in std_logic;
    saxigp5_arcache : in std_logic_vector(3 downto 0);
    saxigp5_arprot : in std_logic_vector(2 downto 0);
    saxigp5_arvalid : in std_logic;
    saxigp5_arready : out std_logic;
    saxigp5_rid : out std_logic_vector(5 downto 0);
    saxigp5_rdata : out std_logic_vector(C_SAXIGP5_DATA_WIDTH-1 downto 0);
    saxigp5_rresp : out std_logic_vector(1 downto 0);
    saxigp5_rlast : out std_logic;
    saxigp5_rvalid : out std_logic;
    saxigp5_rready : in std_logic;
    saxigp5_awqos : in std_logic_vector(3 downto 0);
    saxigp5_arqos : in std_logic_vector(3 downto 0);
    saxigp5_rcount : out std_logic_vector(7 downto 0);
    saxigp5_wcount : out std_logic_vector(7 downto 0);
    saxigp5_racount : out std_logic_vector(3 downto 0);
    saxigp5_wacount : out std_logic_vector(3 downto 0);
-- saxigp6
    saxi_lpd_aclk : in std_logic;
    saxi_lpd_rclk : in std_logic;
    saxi_lpd_wclk : in std_logic;
    saxigp6_aruser : in std_logic;
    saxigp6_awuser : in std_logic;
    saxigp6_awid : in std_logic_vector(5 downto 0);
    saxigp6_awaddr : in std_logic_vector(48 downto 0);
    saxigp6_awlen : in std_logic_vector(7 downto 0);
    saxigp6_awsize : in std_logic_vector(2 downto 0);
    saxigp6_awburst : in std_logic_vector(1 downto 0);
    saxigp6_awlock : in std_logic;
    saxigp6_awcache : in std_logic_vector(3 downto 0);
    saxigp6_awprot : in std_logic_vector(2 downto 0);
    saxigp6_awvalid : in std_logic;
    saxigp6_awready : out std_logic;
    saxigp6_wdata : in std_logic_vector(C_SAXIGP6_DATA_WIDTH-1 downto 0);
    saxigp6_wstrb : in std_logic_vector((C_SAXIGP6_DATA_WIDTH/8) -1  downto 0);
    saxigp6_wlast : in std_logic;
    saxigp6_wvalid : in std_logic;
    saxigp6_wready : out std_logic;
    saxigp6_bid : out std_logic_vector(5 downto 0);
    saxigp6_bresp : out std_logic_vector(1 downto 0);
    saxigp6_bvalid : out std_logic;
    saxigp6_bready : in std_logic;
    saxigp6_arid : in std_logic_vector(5 downto 0);
    saxigp6_araddr : in std_logic_vector(48 downto 0);
    saxigp6_arlen : in std_logic_vector(7 downto 0);
    saxigp6_arsize : in std_logic_vector(2 downto 0);
    saxigp6_arburst : in std_logic_vector(1 downto 0);
    saxigp6_arlock : in std_logic;
    saxigp6_arcache : in std_logic_vector(3 downto 0);
    saxigp6_arprot : in std_logic_vector(2 downto 0);
    saxigp6_arvalid : in std_logic;
    saxigp6_arready : out std_logic;
    saxigp6_rid : out std_logic_vector(5 downto 0);
    saxigp6_rdata : out std_logic_vector(C_SAXIGP6_DATA_WIDTH-1 downto 0);
    saxigp6_rresp : out std_logic_vector(1 downto 0);
    saxigp6_rlast : out std_logic;
    saxigp6_rvalid : out std_logic;
    saxigp6_rready : in std_logic;
    saxigp6_awqos : in std_logic_vector(3 downto 0);
    saxigp6_arqos : in std_logic_vector(3 downto 0);
    saxigp6_rcount : out std_logic_vector(7 downto 0);
    saxigp6_wcount : out std_logic_vector(7 downto 0);
    saxigp6_racount : out std_logic_vector(3 downto 0);
    saxigp6_wacount : out std_logic_vector(3 downto 0);
-- saxiacp
    saxiacp_fpd_aclk : in std_logic;
    saxiacp_awaddr : in std_logic_vector(39 downto 0);
    saxiacp_awid : in std_logic_vector(4 downto 0);
    saxiacp_awlen : in std_logic_vector(7 downto 0);
    saxiacp_awsize : in std_logic_vector(2 downto 0);
    saxiacp_awburst : in std_logic_vector(1 downto 0);
    saxiacp_awlock : in std_logic;
    saxiacp_awcache : in std_logic_vector(3 downto 0);
    saxiacp_awprot : in std_logic_vector(2 downto 0);
    saxiacp_awvalid : in std_logic;
    saxiacp_awready : out std_logic;
    saxiacp_awuser : in std_logic_vector(1 downto 0);
    saxiacp_awqos : in std_logic_vector(3 downto 0);
    saxiacp_wlast : in std_logic;
    saxiacp_wdata : in std_logic_vector(127 downto 0);
    saxiacp_wstrb : in std_logic_vector(15 downto 0);
    saxiacp_wvalid : in std_logic;
    saxiacp_wready : out std_logic;
    saxiacp_bresp : out std_logic_vector(1 downto 0);
    saxiacp_bid : out std_logic_vector(4 downto 0);
    saxiacp_bvalid : out std_logic;
    saxiacp_bready : in std_logic;
    saxiacp_araddr : in std_logic_vector(39 downto 0);
    saxiacp_arid : in std_logic_vector(4 downto 0);
    saxiacp_arlen : in std_logic_vector(7 downto 0);
    saxiacp_arsize : in std_logic_vector(2 downto 0);
    saxiacp_arburst : in std_logic_vector(1 downto 0);
    saxiacp_arlock : in std_logic;
    saxiacp_arcache : in std_logic_vector(3 downto 0);
    saxiacp_arprot : in std_logic_vector(2 downto 0);
    saxiacp_arvalid : in std_logic;
    saxiacp_arready : out std_logic;
    saxiacp_aruser : in std_logic_vector(1 downto 0);
    saxiacp_arqos : in std_logic_vector(3 downto 0);
    saxiacp_rid : out std_logic_vector(4 downto 0);
    saxiacp_rlast : out std_logic;
    saxiacp_rdata : out std_logic_vector(127 downto 0);
    saxiacp_rresp : out std_logic_vector(1 downto 0);
    saxiacp_rvalid : out std_logic;
    saxiacp_rready : in std_logic;
-- sacefpd
    sacefpd_aclk : in std_logic;
    sacefpd_awvalid : in std_logic;
    sacefpd_awready : out std_logic;
    sacefpd_awid : in std_logic_vector(5 downto 0);
    sacefpd_awaddr : in std_logic_vector(43 downto 0);
    sacefpd_awregion : in std_logic_vector(3 downto 0);
    sacefpd_awlen : in std_logic_vector(7 downto 0);
    sacefpd_awsize : in std_logic_vector(2 downto 0);
    sacefpd_awburst : in std_logic_vector(1 downto 0);
    sacefpd_awlock : in std_logic;
    sacefpd_awcache : in std_logic_vector(3 downto 0);
    sacefpd_awprot : in std_logic_vector(2 downto 0);
    sacefpd_awdomain : in std_logic_vector(1 downto 0);
    sacefpd_awsnoop : in std_logic_vector(2 downto 0);
    sacefpd_awbar : in std_logic_vector(1 downto 0);
    sacefpd_awqos : in std_logic_vector(3 downto 0);
    sacefpd_wvalid : in std_logic;
    sacefpd_wready : out std_logic;
    sacefpd_wdata : in std_logic_vector(127 downto 0);
    sacefpd_wstrb : in std_logic_vector(15 downto 0);
    sacefpd_wlast : in std_logic;
    sacefpd_wuser : in std_logic;
    sacefpd_bvalid : out std_logic;
    sacefpd_bready : in std_logic;
    sacefpd_bid : out std_logic_vector(5 downto 0);
    sacefpd_bresp : out std_logic_vector(1 downto 0);
    sacefpd_buser : out std_logic;
    sacefpd_arvalid : in std_logic;
    sacefpd_arready : out std_logic;
    sacefpd_arid : in std_logic_vector(5 downto 0);
    sacefpd_araddr : in std_logic_vector(43 downto 0);
    sacefpd_arregion : in std_logic_vector(3 downto 0);
    sacefpd_arlen : in std_logic_vector(7 downto 0);
    sacefpd_arsize : in std_logic_vector(2 downto 0);
    sacefpd_arburst : in std_logic_vector(1 downto 0);
    sacefpd_arlock : in std_logic;
    sacefpd_arcache : in std_logic_vector(3 downto 0);
    sacefpd_arprot : in std_logic_vector(2 downto 0);
    sacefpd_ardomain : in std_logic_vector(1 downto 0);
    sacefpd_arsnoop : in std_logic_vector(3 downto 0);
    sacefpd_arbar : in std_logic_vector(1 downto 0);
    sacefpd_arqos : in std_logic_vector(3 downto 0);
    sacefpd_rvalid : out std_logic;
    sacefpd_rready : in std_logic;
    sacefpd_rid : out std_logic_vector(5 downto 0);
    sacefpd_rdata : out std_logic_vector(127 downto 0);
    sacefpd_rresp : out std_logic_vector(3 downto 0);
    sacefpd_rlast : out std_logic;
    sacefpd_ruser : out std_logic;
    sacefpd_acvalid : out std_logic;
    sacefpd_acready : in std_logic;
    sacefpd_acaddr : out std_logic_vector(43 downto 0);
    sacefpd_acsnoop : out std_logic_vector(3 downto 0);
    sacefpd_acprot : out std_logic_vector(2 downto 0);
    sacefpd_crvalid : in std_logic;
    sacefpd_crready : out std_logic;
    sacefpd_crresp : in std_logic_vector(4 downto 0);
    sacefpd_cdvalid : in std_logic;
    sacefpd_cdready : out std_logic;
    sacefpd_cddata : in std_logic_vector(127 downto 0);
    sacefpd_cdlast : in std_logic;
    sacefpd_wack : in std_logic;
    sacefpd_rack : in std_logic;


-----------------------------------------------
-- not using anything below this line yet... --
-----------------------------------------------

-- can0
    emio_can0_phy_tx : out std_logic;
    emio_can0_phy_rx : in std_logic;
-- can1
    emio_can1_phy_tx : out std_logic;
    emio_can1_phy_rx : in std_logic;
-- enet0
    emio_enet0_gmii_rx_clk : in std_logic;
    emio_enet0_speed_mode : out std_logic_vector(2 downto 0);
    emio_enet0_gmii_crs : in std_logic;
    emio_enet0_gmii_col : in std_logic;
    emio_enet0_gmii_rxd : in std_logic_vector(7 downto 0);
    emio_enet0_gmii_rx_er : in std_logic;
    emio_enet0_gmii_rx_dv : in std_logic;
    emio_enet0_gmii_tx_clk : in std_logic;
    emio_enet0_gmii_txd : out std_logic_vector(7 downto 0);
    emio_enet0_gmii_tx_en : out std_logic;
    emio_enet0_gmii_tx_er : out std_logic;
    emio_enet0_mdio_mdc : out std_logic;
    emio_enet0_mdio_i : in std_logic;
    emio_enet0_mdio_o : out std_logic;
    emio_enet0_mdio_t : out std_logic;
    emio_enet0_mdio_t_n : out std_logic;
-- enet1
    emio_enet1_gmii_rx_clk : in std_logic;
    emio_enet1_speed_mode : out std_logic_vector(2 downto 0);
    emio_enet1_gmii_crs : in std_logic;
    emio_enet1_gmii_col : in std_logic;
    emio_enet1_gmii_rxd : in std_logic_vector(7 downto 0);
    emio_enet1_gmii_rx_er : in std_logic;
    emio_enet1_gmii_rx_dv : in std_logic;
    emio_enet1_gmii_tx_clk : in std_logic;
    emio_enet1_gmii_txd : out std_logic_vector(7 downto 0);
    emio_enet1_gmii_tx_en : out std_logic;
    emio_enet1_gmii_tx_er : out std_logic;
    emio_enet1_mdio_mdc : out std_logic;
    emio_enet1_mdio_i : in std_logic;
    emio_enet1_mdio_o : out std_logic;
    emio_enet1_mdio_t : out std_logic;
    emio_enet1_mdio_t_n : out std_logic;
-- enet2
    emio_enet2_gmii_rx_clk : in std_logic;
    emio_enet2_speed_mode : out std_logic_vector(2 downto 0);
    emio_enet2_gmii_crs : in std_logic;
    emio_enet2_gmii_col : in std_logic;
    emio_enet2_gmii_rxd : in std_logic_vector(7 downto 0);
    emio_enet2_gmii_rx_er : in std_logic;
    emio_enet2_gmii_rx_dv : in std_logic;
    emio_enet2_gmii_tx_clk : in std_logic;
    emio_enet2_gmii_txd : out std_logic_vector(7 downto 0);
    emio_enet2_gmii_tx_en : out std_logic;
    emio_enet2_gmii_tx_er : out std_logic;
    emio_enet2_mdio_mdc : out std_logic;
    emio_enet2_mdio_i : in std_logic;
    emio_enet2_mdio_o : out std_logic;
    emio_enet2_mdio_t : out std_logic;
    emio_enet2_mdio_t_n : out std_logic;
-- enet3
    emio_enet3_gmii_rx_clk : in std_logic;
    emio_enet3_speed_mode : out std_logic_vector(2 downto 0);
    emio_enet3_gmii_crs : in std_logic;
    emio_enet3_gmii_col : in std_logic;
    emio_enet3_gmii_rxd : in std_logic_vector(7 downto 0);
    emio_enet3_gmii_rx_er : in std_logic;
    emio_enet3_gmii_rx_dv : in std_logic;
    emio_enet3_gmii_tx_clk : in std_logic;
    emio_enet3_gmii_txd : out std_logic_vector(7 downto 0);
    emio_enet3_gmii_tx_en : out std_logic;
    emio_enet3_gmii_tx_er : out std_logic;
    emio_enet3_mdio_mdc : out std_logic;
    emio_enet3_mdio_i : in std_logic;
    emio_enet3_mdio_o : out std_logic;
    emio_enet3_mdio_t : out std_logic;
    emio_enet3_mdio_t_n : out std_logic;
-- fifoif0
    emio_enet0_tx_r_data_rdy : in std_logic;
    emio_enet0_tx_r_rd : out std_logic;
    emio_enet0_tx_r_valid : in std_logic;
    emio_enet0_tx_r_data : in std_logic_vector(7 downto 0);
    emio_enet0_tx_r_sop : in std_logic;
    emio_enet0_tx_r_eop : in std_logic;
    emio_enet0_tx_r_err : in std_logic;
    emio_enet0_tx_r_underflow : in std_logic;
    emio_enet0_tx_r_flushed : in std_logic;
    emio_enet0_tx_r_control : in std_logic;
    emio_enet0_dma_tx_end_tog : out std_logic;
    emio_enet0_dma_tx_status_tog : in std_logic;
    emio_enet0_tx_r_status : out std_logic_vector(3 downto 0);
    emio_enet0_rx_w_wr : out std_logic;
    emio_enet0_rx_w_data : out std_logic_vector(7 downto 0);
    emio_enet0_rx_w_sop : out std_logic;
    emio_enet0_rx_w_eop : out std_logic;
    emio_enet0_rx_w_status : out std_logic_vector(44 downto 0);
    emio_enet0_rx_w_err : out std_logic;
    emio_enet0_rx_w_overflow : in std_logic;
    emio_enet0_signal_detect : in std_logic;
    emio_enet0_rx_w_flush : out std_logic;
    emio_enet0_tx_r_fixed_lat : out std_logic;
-- fifoif1
    emio_enet1_tx_r_data_rdy : in std_logic;
    emio_enet1_tx_r_rd : out std_logic;
    emio_enet1_tx_r_valid : in std_logic;
    emio_enet1_tx_r_data : in std_logic_vector(7 downto 0);
    emio_enet1_tx_r_sop : in std_logic;
    emio_enet1_tx_r_eop : in std_logic;
    emio_enet1_tx_r_err : in std_logic;
    emio_enet1_tx_r_underflow : in std_logic;
    emio_enet1_tx_r_flushed : in std_logic;
    emio_enet1_tx_r_control : in std_logic;
    emio_enet1_dma_tx_end_tog : out std_logic;
    emio_enet1_dma_tx_status_tog : in std_logic;
    emio_enet1_tx_r_status : out std_logic_vector(3 downto 0);
    emio_enet1_rx_w_wr : out std_logic;
    emio_enet1_rx_w_data : out std_logic_vector(7 downto 0);
    emio_enet1_rx_w_sop : out std_logic;
    emio_enet1_rx_w_eop : out std_logic;
    emio_enet1_rx_w_status : out std_logic_vector(44 downto 0);
    emio_enet1_rx_w_err : out std_logic;
    emio_enet1_rx_w_overflow : in std_logic;
    emio_enet1_signal_detect : in std_logic;
    emio_enet1_rx_w_flush : out std_logic;
    emio_enet1_tx_r_fixed_lat : out std_logic;
-- fifoif2
    emio_enet2_tx_r_data_rdy : in std_logic;
    emio_enet2_tx_r_rd : out std_logic;
    emio_enet2_tx_r_valid : in std_logic;
    emio_enet2_tx_r_data : in std_logic_vector(7 downto 0);
    emio_enet2_tx_r_sop : in std_logic;
    emio_enet2_tx_r_eop : in std_logic;
    emio_enet2_tx_r_err : in std_logic;
    emio_enet2_tx_r_underflow : in std_logic;
    emio_enet2_tx_r_flushed : in std_logic;
    emio_enet2_tx_r_control : in std_logic;
    emio_enet2_dma_tx_end_tog : out std_logic;
    emio_enet2_dma_tx_status_tog : in std_logic;
    emio_enet2_tx_r_status : out std_logic_vector(3 downto 0);
    emio_enet2_rx_w_wr : out std_logic;
    emio_enet2_rx_w_data : out std_logic_vector(7 downto 0);
    emio_enet2_rx_w_sop : out std_logic;
    emio_enet2_rx_w_eop : out std_logic;
    emio_enet2_rx_w_status : out std_logic_vector(44 downto 0);
    emio_enet2_rx_w_err : out std_logic;
    emio_enet2_rx_w_overflow : in std_logic;
    emio_enet2_signal_detect : in std_logic;
    emio_enet2_rx_w_flush : out std_logic;
    emio_enet2_tx_r_fixed_lat : out std_logic;
-- fifoif3
    emio_enet3_tx_r_data_rdy : in std_logic;
    emio_enet3_tx_r_rd : out std_logic;
    emio_enet3_tx_r_valid : in std_logic;
    emio_enet3_tx_r_data : in std_logic_vector(7 downto 0);
    emio_enet3_tx_r_sop : in std_logic;
    emio_enet3_tx_r_eop : in std_logic;
    emio_enet3_tx_r_err : in std_logic;
    emio_enet3_tx_r_underflow : in std_logic;
    emio_enet3_tx_r_flushed : in std_logic;
    emio_enet3_tx_r_control : in std_logic;
    emio_enet3_dma_tx_end_tog : out std_logic;
    emio_enet3_dma_tx_status_tog : in std_logic;
    emio_enet3_tx_r_status : out std_logic_vector(3 downto 0);
    emio_enet3_rx_w_wr : out std_logic;
    emio_enet3_rx_w_data : out std_logic_vector(7 downto 0);
    emio_enet3_rx_w_sop : out std_logic;
    emio_enet3_rx_w_eop : out std_logic;
    emio_enet3_rx_w_status : out std_logic_vector(44 downto 0);
    emio_enet3_rx_w_err : out std_logic;
    emio_enet3_rx_w_overflow : in std_logic;
    emio_enet3_signal_detect : in std_logic;
    emio_enet3_rx_w_flush : out std_logic;
    emio_enet3_tx_r_fixed_lat : out std_logic;
-- gem0_fmio
--    fmio_gem0_fifo_tx_clk_from_pl : in std_logic;
--    fmio_gem0_fifo_rx_clk_from_pl : in std_logic;
    fmio_gem0_fifo_tx_clk_to_pl_bufg : out std_logic;
    fmio_gem0_fifo_rx_clk_to_pl_bufg : out std_logic;
-- gem1_fmio
--    fmio_gem1_fifo_tx_clk_from_pl : in std_logic;
--    fmio_gem1_fifo_rx_clk_from_pl : in std_logic;
    fmio_gem1_fifo_tx_clk_to_pl_bufg : out std_logic;
    fmio_gem1_fifo_rx_clk_to_pl_bufg : out std_logic;
-- gem2_fmio
--    fmio_gem2_fifo_tx_clk_from_pl : in std_logic;
--    fmio_gem2_fifo_rx_clk_from_pl : in std_logic;
    fmio_gem2_fifo_tx_clk_to_pl_bufg : out std_logic;
    fmio_gem2_fifo_rx_clk_to_pl_bufg : out std_logic;
-- gem3_fmio
--    fmio_gem3_fifo_tx_clk_from_pl : in std_logic;
--    fmio_gem3_fifo_rx_clk_from_pl : in std_logic;
    fmio_gem3_fifo_tx_clk_to_pl_bufg : out std_logic;
    fmio_gem3_fifo_rx_clk_to_pl_bufg : out std_logic;
-- gem0_1588
     emio_enet0_tx_sof : out std_logic;
     emio_enet0_sync_frame_tx : out std_logic;
     emio_enet0_delay_req_tx : out std_logic;
     emio_enet0_pdelay_req_tx : out std_logic;
     emio_enet0_pdelay_resp_tx : out std_logic;
     emio_enet0_rx_sof : out std_logic;
     emio_enet0_sync_frame_rx : out std_logic;
     emio_enet0_delay_req_rx : out std_logic;
     emio_enet0_pdelay_req_rx : out std_logic;
     emio_enet0_pdelay_resp_rx : out std_logic;
     emio_enet0_tsu_inc_ctrl : in std_logic_vector(1 downto 0);
     emio_enet0_tsu_timer_cmp_val : out std_logic;
--gem1_1588
     emio_enet1_tx_sof : out std_logic;
     emio_enet1_sync_frame_tx : out std_logic;
     emio_enet1_delay_req_tx : out std_logic;
     emio_enet1_pdelay_req_tx : out std_logic;
     emio_enet1_pdelay_resp_tx : out std_logic;
     emio_enet1_rx_sof : out std_logic;
     emio_enet1_sync_frame_rx : out std_logic;
     emio_enet1_delay_req_rx : out std_logic;
     emio_enet1_pdelay_req_rx : out std_logic;
     emio_enet1_pdelay_resp_rx : out std_logic;
     emio_enet1_tsu_inc_ctrl : in std_logic_vector(1 downto 0);
     emio_enet1_tsu_timer_cmp_val : out std_logic;
--gem2_1588
     emio_enet2_tx_sof : out std_logic;
     emio_enet2_sync_frame_tx : out std_logic;
     emio_enet2_delay_req_tx : out std_logic;
     emio_enet2_pdelay_req_tx : out std_logic;
     emio_enet2_pdelay_resp_tx : out std_logic;
     emio_enet2_rx_sof : out std_logic;
     emio_enet2_sync_frame_rx : out std_logic;
     emio_enet2_delay_req_rx : out std_logic;
     emio_enet2_pdelay_req_rx : out std_logic;
     emio_enet2_pdelay_resp_rx : out std_logic;
     emio_enet2_tsu_inc_ctrl : in std_logic_vector(1 downto 0);
     emio_enet2_tsu_timer_cmp_val : out std_logic;
--gem3_1588
     emio_enet3_tx_sof : out std_logic;
     emio_enet3_sync_frame_tx : out std_logic;
     emio_enet3_delay_req_tx : out std_logic;
     emio_enet3_pdelay_req_tx : out std_logic;
     emio_enet3_pdelay_resp_tx : out std_logic;
     emio_enet3_rx_sof : out std_logic;
     emio_enet3_sync_frame_rx : out std_logic;
     emio_enet3_delay_req_rx : out std_logic;
     emio_enet3_pdelay_req_rx : out std_logic;
     emio_enet3_pdelay_resp_rx : out std_logic;
     emio_enet3_tsu_inc_ctrl : in std_logic_vector(1 downto 0);
     emio_enet3_tsu_timer_cmp_val : out std_logic;
-- gem_tsu
    fmio_gem_tsu_clk_from_pl : in std_logic;
    fmio_gem_tsu_clk_to_pl_bufg : out std_logic;
    emio_enet_tsu_clk : in std_logic;
    emio_enet0_enet_tsu_timer_cnt : out std_logic_vector(93 downto 0);
-- gem_misc
    emio_enet0_ext_int_in : in std_logic;
    emio_enet1_ext_int_in : in std_logic;
    emio_enet2_ext_int_in : in std_logic;
    emio_enet3_ext_int_in : in std_logic;
    emio_enet0_dma_bus_width : out std_logic_vector(1 downto 0);
    emio_enet1_dma_bus_width : out std_logic_vector(1 downto 0);
    emio_enet2_dma_bus_width : out std_logic_vector(1 downto 0);
    emio_enet3_dma_bus_width : out std_logic_vector(1 downto 0);
-- gpio
    emio_gpio_i : in std_logic_vector((C_EMIO_GPIO_WIDTH -1) downto 0);
    emio_gpio_o : out std_logic_vector((C_EMIO_GPIO_WIDTH -1) downto 0);
    emio_gpio_t : out std_logic_vector((C_EMIO_GPIO_WIDTH -1) downto 0);
    emio_gpio_t_n : out std_logic_vector((C_EMIO_GPIO_WIDTH -1) downto 0);
-- i2c0
    emio_i2c0_scl_i : in std_logic;
    emio_i2c0_scl_o : out std_logic;
    emio_i2c0_scl_t_n : out std_logic;
    emio_i2c0_scl_t : out std_logic;
    emio_i2c0_sda_i : in std_logic;
    emio_i2c0_sda_o : out std_logic;
    emio_i2c0_sda_t_n : out std_logic;
    emio_i2c0_sda_t : out std_logic;
-- i2c1
    emio_i2c1_scl_i : in std_logic;
    emio_i2c1_scl_o : out std_logic;
    emio_i2c1_scl_t : out std_logic;
    emio_i2c1_scl_t_n : out std_logic;
    emio_i2c1_sda_i : in std_logic;
    emio_i2c1_sda_o : out std_logic;
    emio_i2c1_sda_t : out std_logic;
    emio_i2c1_sda_t_n : out std_logic;
-- uart0
    emio_uart0_txd : out std_logic;
    emio_uart0_rxd : in std_logic;
    emio_uart0_ctsn : in std_logic;
    emio_uart0_rtsn : out std_logic;
    emio_uart0_dsrn : in std_logic;
    emio_uart0_dcdn : in std_logic;
    emio_uart0_rin : in std_logic;
    emio_uart0_dtrn : out std_logic;
-- uart1
    emio_uart1_txd : out std_logic;
    emio_uart1_rxd : in std_logic;
    emio_uart1_ctsn : in std_logic;
    emio_uart1_rtsn : out std_logic;
    emio_uart1_dsrn : in std_logic;
    emio_uart1_dcdn : in std_logic;
    emio_uart1_rin : in std_logic;
    emio_uart1_dtrn : out std_logic;
-- sdio0
    emio_sdio0_clkout : out std_logic;
    emio_sdio0_fb_clk_in : in std_logic;
    emio_sdio0_cmdout : out std_logic;
    emio_sdio0_cmdin : in std_logic;
    emio_sdio0_cmdena : out std_logic;
    emio_sdio0_datain : in std_logic_vector(C_SD0_INTERNAL_BUS_WIDTH-1 downto 0);
    emio_sdio0_dataout : out std_logic_vector(C_SD0_INTERNAL_BUS_WIDTH-1 downto 0);
    emio_sdio0_dataena : out std_logic_vector(C_SD0_INTERNAL_BUS_WIDTH-1 downto 0);
    emio_sdio0_cd_n : in std_logic;
    emio_sdio0_wp : in std_logic;
    emio_sdio0_ledcontrol : out std_logic;
    emio_sdio0_buspower : out std_logic;
    emio_sdio0_bus_volt : out std_logic_vector(2 downto 0);
-- sdio1
    emio_sdio1_clkout : out std_logic;
    emio_sdio1_fb_clk_in : in std_logic;
    emio_sdio1_cmdout : out std_logic;
    emio_sdio1_cmdin : in std_logic;
    emio_sdio1_cmdena : out std_logic;
    emio_sdio1_datain : in std_logic_vector(C_SD1_INTERNAL_BUS_WIDTH-1 downto 0);
    emio_sdio1_dataout : out std_logic_vector(C_SD1_INTERNAL_BUS_WIDTH-1 downto 0);
    emio_sdio1_dataena : out std_logic_vector(C_SD1_INTERNAL_BUS_WIDTH-1 downto 0);
    emio_sdio1_cd_n : in std_logic;
    emio_sdio1_wp : in std_logic;
    emio_sdio1_ledcontrol : out std_logic;
    emio_sdio1_buspower : out std_logic;
    emio_sdio1_bus_volt : out std_logic_vector(2 downto 0);
-- spi0
    emio_spi0_sclk_i : in std_logic;
    emio_spi0_sclk_o : out std_logic;
    emio_spi0_sclk_t : out std_logic;
    emio_spi0_sclk_t_n : out std_logic;
    emio_spi0_m_i : in std_logic;
    emio_spi0_m_o : out std_logic;
    emio_spi0_mo_t : out std_logic;
    emio_spi0_mo_t_n : out std_logic;
    emio_spi0_s_i : in std_logic;
    emio_spi0_s_o : out std_logic;
    emio_spi0_so_t : out std_logic;
    emio_spi0_so_t_n : out std_logic;
    emio_spi0_ss_i_n : in std_logic;
    emio_spi0_ss_o_n : out std_logic;
    emio_spi0_ss1_o_n : out std_logic;
    emio_spi0_ss2_o_n : out std_logic;
    emio_spi0_ss_n_t : out std_logic;
    emio_spi0_ss_n_t_n : out std_logic;
-- spi1
    emio_spi1_sclk_i : in std_logic;
    emio_spi1_sclk_o : out std_logic;
    emio_spi1_sclk_t : out std_logic;
    emio_spi1_sclk_t_n : out std_logic;
    emio_spi1_m_i : in std_logic;
    emio_spi1_m_o : out std_logic;
    emio_spi1_mo_t : out std_logic;
    emio_spi1_mo_t_n : out std_logic;
    emio_spi1_s_i : in std_logic;
    emio_spi1_s_o : out std_logic;
    emio_spi1_so_t : out std_logic;
    emio_spi1_so_t_n : out std_logic;
    emio_spi1_ss_i_n : in std_logic;
    emio_spi1_ss_o_n : out std_logic;
    emio_spi1_ss1_o_n : out std_logic;
    emio_spi1_ss2_o_n : out std_logic;
    emio_spi1_ss_n_t : out std_logic;
    emio_spi1_ss_n_t_n : out std_logic;
-- trace
    pl_ps_trace_clk : in std_logic;
    ps_pl_tracectl : out std_logic;
    ps_pl_tracedata : out std_logic_vector(C_TRACE_DATA_WIDTH-1 downto 0);
    trace_clk_out : out std_logic;
-- ttc0
    emio_ttc0_wave_o : out std_logic_vector(2 downto 0);
    emio_ttc0_clk_i : in std_logic_vector(2 downto 0);
-- ttc1
    emio_ttc1_wave_o : out std_logic_vector(2 downto 0);
    emio_ttc1_clk_i : in std_logic_vector(2 downto 0);
-- ttc2
    emio_ttc2_wave_o : out std_logic_vector(2 downto 0);
    emio_ttc2_clk_i : in std_logic_vector(2 downto 0);
-- ttc3
    emio_ttc3_wave_o : out std_logic_vector(2 downto 0);
    emio_ttc3_clk_i : in std_logic_vector(2 downto 0);
-- wdt0
    emio_wdt0_clk_i : in std_logic;
    emio_wdt0_rst_o : out std_logic;
-- wdt1
    emio_wdt1_clk_i : in std_logic;
    emio_wdt1_rst_o : out std_logic;
-- usb3
    emio_hub_port_overcrnt_usb3_0 : in std_logic;
    emio_hub_port_overcrnt_usb3_1 : in std_logic;
    emio_hub_port_overcrnt_usb2_0 : in std_logic;
    emio_hub_port_overcrnt_usb2_1 : in std_logic;
    emio_u2dsport_vbus_ctrl_usb3_0 : out std_logic;
    emio_u2dsport_vbus_ctrl_usb3_1 : out std_logic;
    emio_u3dsport_vbus_ctrl_usb3_0 : out std_logic;
    emio_u3dsport_vbus_ctrl_usb3_1 : out std_logic;
--adma
    adma_fci_clk : in std_logic_vector(7 downto 0);
    pl2adma_cvld : in std_logic_vector(7 downto 0);
    pl2adma_tack : in std_logic_vector(7 downto 0);
    adma2pl_cack : out std_logic_vector(7 downto 0);
    adma2pl_tvld : out std_logic_vector(7 downto 0);
--gdma
    perif_gdma_clk : in std_logic_vector(7 downto 0);
    perif_gdma_cvld : in std_logic_vector(7 downto 0);
    perif_gdma_tack : in std_logic_vector(7 downto 0);
    gdma_perif_cack : out std_logic_vector(7 downto 0);
    gdma_perif_tvld : out std_logic_vector(7 downto 0);
-- clk
    pl_clock_stop : in std_logic_vector(3 downto 0);
    pll_aux_refclk_lpd : in std_logic_vector(1 downto 0);
    pll_aux_refclk_fpd : in std_logic_vector(2 downto 0);
-- audio
    dp_s_axis_audio_tdata : in std_logic_vector(31 downto 0);
    dp_s_axis_audio_tid : in std_logic;
    dp_s_axis_audio_tvalid : in std_logic;
    dp_s_axis_audio_tready : out std_logic;
    dp_m_axis_mixed_audio_tdata : out std_logic_vector(31 downto 0);
    dp_m_axis_mixed_audio_tid : out std_logic;
    dp_m_axis_mixed_audio_tvalid : out std_logic;
    dp_m_axis_mixed_audio_tready : in std_logic;
    dp_s_axis_audio_clk : in std_logic;
-- video
    dp_live_video_in_vsync : in std_logic;
    dp_live_video_in_hsync : in std_logic;
    dp_live_video_in_de : in std_logic;
    dp_live_video_in_pixel1 : in std_logic_vector(35 downto 0);
    dp_video_in_clk : in std_logic;
    dp_video_out_hsync : out std_logic;
    dp_video_out_vsync : out std_logic;
    dp_video_out_pixel1 : out std_logic_vector(35 downto 0);
    dp_aux_data_in : in std_logic;
    dp_aux_data_out : out std_logic;
    dp_aux_data_oe_n : out std_logic;
    dp_live_gfx_alpha_in : in std_logic_vector(7 downto 0);
    dp_live_gfx_pixel1_in : in std_logic_vector(35 downto 0);
    dp_hot_plug_detect : in std_logic;
    dp_external_custom_event1 : in std_logic;
    dp_external_custom_event2 : in std_logic;
    dp_external_vsync_event : in std_logic;
    dp_live_video_de_out : out std_logic;
-- event_apu
    pl_ps_eventi : in std_logic;
    ps_pl_evento : out std_logic;
    ps_pl_standbywfe : out std_logic_vector(3 downto 0);
    ps_pl_standbywfi : out std_logic_vector(3 downto 0);
    pl_ps_apugic_irq : in std_logic_vector(3 downto 0);
    pl_ps_apugic_fiq : in std_logic_vector(3 downto 0);
-- event_rpu
    rpu_eventi0 : in std_logic;
    rpu_eventi1 : in std_logic;
    rpu_evento0 : out std_logic;
    rpu_evento1 : out std_logic;
    nfiq0_lpd_rpu : in std_logic;
    nfiq1_lpd_rpu : in std_logic;
    nirq0_lpd_rpu : in std_logic;
    nirq1_lpd_rpu : in std_logic;
-- ipi
    irq_ipi_pl_0 : out std_logic;
    irq_ipi_pl_1 : out std_logic;
    irq_ipi_pl_2 : out std_logic;
    irq_ipi_pl_3 : out std_logic;
-- stm
    stm_event : in std_logic_vector(59 downto 0);
-- ftm
    pl_ps_trigack_0 : in std_logic;
    pl_ps_trigack_1 : in std_logic;
    pl_ps_trigack_2 : in std_logic;
    pl_ps_trigack_3 : in std_logic;
    pl_ps_trigger_0 : in std_logic;
    pl_ps_trigger_1 : in std_logic;
    pl_ps_trigger_2 : in std_logic;
    pl_ps_trigger_3 : in std_logic;
    ps_pl_trigack_0 : out std_logic;
    ps_pl_trigack_1 : out std_logic;
    ps_pl_trigack_2 : out std_logic;
    ps_pl_trigack_3 : out std_logic;
    ps_pl_trigger_0 : out std_logic;
    ps_pl_trigger_1 : out std_logic;
    ps_pl_trigger_2 : out std_logic;
    ps_pl_trigger_3 : out std_logic;
    ftm_gpo : out std_logic_vector(31 downto 0);
    ftm_gpi : in std_logic_vector(31 downto 0);
-- irq
    pl_ps_irq0 : in std_logic_vector((C_NUM_F2P_0_INTR_INPUTS-1) downto 0);
    pl_ps_irq1 : in std_logic_vector((C_NUM_F2P_1_INTR_INPUTS-1) downto 0);
--    ps_pl_irq_lpd : out std_logic_vector(99 downto 0);
--    ps_pl_irq_fpd : out std_logic_vector(63 downto 0);

--resets using gpio

    pl_resetn0 : out std_logic;
    pl_resetn1 : out std_logic;
    pl_resetn2 : out std_logic;
    pl_resetn3 : out std_logic;

    ps_pl_irq_can0 : out std_logic;
    ps_pl_irq_can1 : out std_logic;
    ps_pl_irq_enet0 : out std_logic;
    ps_pl_irq_enet1 : out std_logic;
    ps_pl_irq_enet2 : out std_logic;
    ps_pl_irq_enet3 : out std_logic;
    ps_pl_irq_enet0_wake : out std_logic;
    ps_pl_irq_enet1_wake : out std_logic;
    ps_pl_irq_enet2_wake : out std_logic;
    ps_pl_irq_enet3_wake : out std_logic;
    ps_pl_irq_gpio : out std_logic;
    ps_pl_irq_i2c0 : out std_logic;
    ps_pl_irq_i2c1 : out std_logic;
    ps_pl_irq_uart0 : out std_logic;
    ps_pl_irq_uart1 : out std_logic;
    ps_pl_irq_sdio0 : out std_logic;
    ps_pl_irq_sdio1 : out std_logic;
    ps_pl_irq_sdio0_wake : out std_logic;
    ps_pl_irq_sdio1_wake : out std_logic;
    ps_pl_irq_spi0 : out std_logic;
    ps_pl_irq_spi1 : out std_logic;
    ps_pl_irq_qspi : out std_logic;
    ps_pl_irq_ttc0_0 : out std_logic;
    ps_pl_irq_ttc0_1 : out std_logic;
    ps_pl_irq_ttc0_2 : out std_logic;
    ps_pl_irq_ttc1_0 : out std_logic;
    ps_pl_irq_ttc1_1 : out std_logic;
    ps_pl_irq_ttc1_2 : out std_logic;
    ps_pl_irq_ttc2_0 : out std_logic;
    ps_pl_irq_ttc2_1 : out std_logic;
    ps_pl_irq_ttc2_2 : out std_logic;
    ps_pl_irq_ttc3_0 : out std_logic;
    ps_pl_irq_ttc3_1 : out std_logic;
    ps_pl_irq_ttc3_2 : out std_logic;
    ps_pl_irq_csu_pmu_wdt : out std_logic;
    ps_pl_irq_lp_wdt : out std_logic;
    ps_pl_irq_usb3_0_endpoint : out std_logic_vector(3 downto 0);
    ps_pl_irq_usb3_0_otg : out std_logic;
    ps_pl_irq_usb3_1_endpoint : out std_logic_vector(3 downto 0);
    ps_pl_irq_usb3_1_otg : out std_logic;
    ps_pl_irq_adma_chan : out std_logic_vector(7 downto 0);
    ps_pl_irq_usb3_0_pmu_wakeup : out std_logic_vector(1 downto 0);
    ps_pl_irq_gdma_chan : out std_logic_vector(7 downto 0);
    ps_pl_irq_csu : out std_logic;
    ps_pl_irq_csu_dma : out std_logic;
    ps_pl_irq_efuse : out std_logic;
    ps_pl_irq_xmpu_lpd : out std_logic;
    ps_pl_irq_ddr_ss : out std_logic;
    ps_pl_irq_nand : out std_logic;
    ps_pl_irq_fp_wdt : out std_logic;
    ps_pl_irq_pcie_msi : out std_logic_vector(1 downto 0);
    ps_pl_irq_pcie_legacy : out std_logic;
    ps_pl_irq_pcie_dma : out std_logic;
    ps_pl_irq_pcie_msc : out std_logic;
    ps_pl_irq_dport : out std_logic;
    ps_pl_irq_fpd_apb_int : out std_logic;
    ps_pl_irq_fpd_atb_error : out std_logic;
    ps_pl_irq_dpdma : out std_logic;
    ps_pl_irq_apm_fpd : out std_logic;
    ps_pl_irq_gpu : out std_logic;
    ps_pl_irq_sata : out std_logic;
    ps_pl_irq_xmpu_fpd : out std_logic;
    ps_pl_irq_apu_cpumnt : out std_logic_vector(3 downto 0);
    ps_pl_irq_apu_cti : out std_logic_vector(3 downto 0);
    ps_pl_irq_apu_pmu : out std_logic_vector(3 downto 0);
    ps_pl_irq_apu_comm : out std_logic_vector(3 downto 0);
    ps_pl_irq_apu_l2err : out std_logic;
    ps_pl_irq_apu_exterr : out std_logic;
    ps_pl_irq_apu_regs : out std_logic;
    ps_pl_irq_intf_ppd_cci : out std_logic;
    ps_pl_irq_intf_fpd_smmu : out std_logic;
    ps_pl_irq_atb_err_lpd : out std_logic;
    ps_pl_irq_aib_axi : out std_logic;
    ps_pl_irq_ams : out std_logic;
    ps_pl_irq_lpd_apm : out std_logic;
    ps_pl_irq_rtc_alaram : out std_logic;
    ps_pl_irq_rtc_seconds : out std_logic;
    ps_pl_irq_clkmon : out std_logic;
    ps_pl_irq_ipi_channel0 : out std_logic;
    ps_pl_irq_ipi_channel1 : out std_logic;
    ps_pl_irq_ipi_channel2 : out std_logic;
    ps_pl_irq_ipi_channel7 : out std_logic;
    ps_pl_irq_ipi_channel8 : out std_logic;
    ps_pl_irq_ipi_channel9 : out std_logic;
    ps_pl_irq_ipi_channel10 : out std_logic;
    ps_pl_irq_rpu_pm : out std_logic_vector(1 downto 0);
    ps_pl_irq_ocm_error : out std_logic;
    ps_pl_irq_lpd_apb_intr : out std_logic;
    ps_pl_irq_r5_core0_ecc_error : out std_logic;
    ps_pl_irq_r5_core1_ecc_error : out std_logic;


-- rtc
    osc_rtc_clk : out std_logic;
-- pmu
    pl_pmu_gpi : in std_logic_vector(31 downto 0);
    pmu_pl_gpo : out std_logic_vector(31 downto 0);
    aib_pmu_afifm_fpd_ack : in std_logic;
    aib_pmu_afifm_lpd_ack : in std_logic;
    pmu_aib_afifm_fpd_req : out std_logic;
    pmu_aib_afifm_lpd_req : out std_logic;
    pmu_error_to_pl : out std_logic_vector(46 downto 0);
    pmu_error_from_pl : in std_logic_vector(3 downto 0);
-- misc
    ddrc_ext_refresh_rank0_req : in std_logic;
    ddrc_ext_refresh_rank1_req : in std_logic;
    ddrc_refresh_pl_clk : in std_logic;
    pl_acpinact : in std_logic;

--For Clock buffering
--FCLK
    pl_clk3 : out std_logic;
    pl_clk2 : out std_logic;
    pl_clk1 : out std_logic;
    pl_clk0 : out std_logic;

---------------------------
-- ACE interface allotment
--------------------------
    sacefpd_awuser : in std_logic_vector(15 downto 0);
    sacefpd_aruser : in std_logic_vector(15 downto 0);

--Debug and Test signals
    test_adc_clk : in std_logic_vector(3 downto 0);
    test_adc_in : in std_logic_vector(31 downto 0);
    test_adc2_in : in std_logic_vector(31 downto 0);
    test_db : out std_logic_vector(15 downto 0);
    test_adc_out : out std_logic_vector(19 downto 0);
    test_ams_osc : out std_logic_vector(7 downto 0);
    test_mon_data : out std_logic_vector(15 downto 0);
    test_dclk : in std_logic;
    test_den : in std_logic;
    test_dwe : in std_logic;
    test_daddr : in std_logic_vector(7 downto 0);
    test_di : in std_logic_vector(15 downto 0);
    test_drdy : out std_logic;
    test_do : out std_logic_vector(15 downto 0);
    test_convst : in std_logic;
    pstp_pl_clk : in std_logic_vector(3 downto 0);
    pstp_pl_in : in std_logic_vector(31 downto 0);
    pstp_pl_out : out std_logic_vector(31 downto 0);
    pstp_pl_ts : in std_logic_vector(31 downto 0);
    fmio_test_gem_scanmux_1 : in std_logic;
    fmio_test_gem_scanmux_2 : in std_logic;
    test_char_mode_fpd_n : in std_logic;
    test_char_mode_lpd_n : in std_logic;
    fmio_test_io_char_scan_clock : in std_logic;
    fmio_test_io_char_scanenable : in std_logic;
    fmio_test_io_char_scan_in : in std_logic;
    fmio_test_io_char_scan_out : out std_logic;
    fmio_test_io_char_scan_reset_n : in std_logic;
    fmio_char_afifslpd_test_select_n : in std_logic;
    fmio_char_afifslpd_test_input : in std_logic;
    fmio_char_afifslpd_test_output : out std_logic;
    fmio_char_afifsfpd_test_select_n : in std_logic;
    fmio_char_afifsfpd_test_input : in std_logic;
    fmio_char_afifsfpd_test_output : out std_logic;
    io_char_audio_in_test_data : in std_logic;
    io_char_audio_mux_sel_n : in std_logic;
    io_char_video_in_test_data : in std_logic;
    io_char_video_mux_sel_n : in std_logic;
    io_char_video_out_test_data : out std_logic;
    io_char_audio_out_test_data : out std_logic;
    fmio_test_qspi_scanmux_1_n : in std_logic;
    fmio_test_sdio_scanmux_1 : in std_logic;
    fmio_test_sdio_scanmux_2 : in std_logic;
    fmio_sd0_dll_test_in_n : in std_logic_vector(3 downto 0);
    fmio_sd0_dll_test_out : out std_logic_vector(7 downto 0);
    fmio_sd1_dll_test_in_n : in std_logic_vector(3 downto 0);
    fmio_sd1_dll_test_out : out std_logic_vector(7 downto 0);
    test_pl_scan_chopper_si : in std_logic;
    test_pl_scan_chopper_so : out std_logic;
    test_pl_scan_chopper_trig : in std_logic;
    test_pl_scan_clk0 : in std_logic;
    test_pl_scan_clk1 : in std_logic;
    test_pl_scan_edt_clk : in std_logic;
    test_pl_scan_edt_in_apu : in std_logic;
    test_pl_scan_edt_in_cpu : in std_logic;
    test_pl_scan_edt_in_ddr : in std_logic_vector(3 downto 0);
    test_pl_scan_edt_in_fp : in std_logic_vector(9 downto 0);
    test_pl_scan_edt_in_gpu : in std_logic_vector(3 downto 0);
    test_pl_scan_edt_in_lp : in std_logic_vector(8 downto 0);
    test_pl_scan_edt_in_usb3 : in std_logic_vector(1 downto 0);
    test_pl_scan_edt_out_apu : out std_logic;
    test_pl_scan_edt_out_cpu0 : out std_logic;
    test_pl_scan_edt_out_cpu1 : out std_logic;
    test_pl_scan_edt_out_cpu2 : out std_logic;
    test_pl_scan_edt_out_cpu3 : out std_logic;
    test_pl_scan_edt_out_ddr : out std_logic_vector(3 downto 0);
    test_pl_scan_edt_out_fp : out std_logic_vector(9 downto 0);
    test_pl_scan_edt_out_gpu : out std_logic_vector(3 downto 0);
    test_pl_scan_edt_out_lp : out std_logic_vector(8 downto 0);
    test_pl_scan_edt_out_usb3 : out std_logic_vector(1 downto 0);
    test_pl_scan_edt_update : in std_logic;
    test_pl_scan_reset_n : in std_logic;
    test_pl_scanenable : in std_logic;
    test_pl_scan_pll_reset : in std_logic;
    test_pl_scan_spare_in0 : in std_logic;
    test_pl_scan_spare_in1 : in std_logic;
    test_pl_scan_spare_out0 : out std_logic;
    test_pl_scan_spare_out1 : out std_logic;
    test_pl_scan_wrap_clk : in std_logic;
    test_pl_scan_wrap_ishift : in std_logic;
    test_pl_scan_wrap_oshift : in std_logic;
    test_pl_scan_slcr_config_clk : in std_logic;
    test_pl_scan_slcr_config_rstn : in std_logic;
    test_pl_scan_slcr_config_si : in std_logic;
    test_pl_scan_spare_in2 : in std_logic;
    test_pl_scanenable_slcr_en : in std_logic;
    test_pl_pll_lock_out : out std_logic_vector(4 downto 0);
    test_pl_scan_slcr_config_so : out std_logic;
    tst_rtc_calibreg_in : in std_logic_vector(20 downto 0);
    tst_rtc_calibreg_out : out std_logic_vector(20 downto 0);
    tst_rtc_calibreg_we : in std_logic;
    tst_rtc_clk : in std_logic;
    tst_rtc_osc_clk_out : out std_logic;
    tst_rtc_sec_counter_out : out std_logic_vector(31 downto 0);
    tst_rtc_seconds_raw_int : out std_logic;
    tst_rtc_testclock_select_n : in std_logic;
    tst_rtc_tick_counter_out : out std_logic_vector(15 downto 0);
    tst_rtc_timesetreg_in : in std_logic_vector(31 downto 0);
    tst_rtc_timesetreg_out : out std_logic_vector(31 downto 0);
    tst_rtc_disable_bat_op : in std_logic;
    tst_rtc_osc_cntrl_in : in std_logic_vector(3 downto 0);
    tst_rtc_osc_cntrl_out : out std_logic_vector(3 downto 0);
    tst_rtc_osc_cntrl_we : in std_logic;
    tst_rtc_sec_reload : in std_logic;
    tst_rtc_timesetreg_we : in std_logic;
    tst_rtc_testmode_n : in std_logic;
    test_usb0_funcmux_0_n : in std_logic;
    test_usb1_funcmux_0_n : in std_logic;
    test_usb0_scanmux_0_n : in std_logic;
    test_usb1_scanmux_0_n : in std_logic;
    lpd_pll_test_out : out std_logic_vector(31 downto 0);
    pl_lpd_pll_test_ck_sel_n : in std_logic_vector(2 downto 0);
    pl_lpd_pll_test_fract_clk_sel_n : in std_logic;
    pl_lpd_pll_test_fract_en_n : in std_logic;
    pl_lpd_pll_test_mux_sel : in std_logic;
    pl_lpd_pll_test_sel : in std_logic_vector(3 downto 0);
    fpd_pll_test_out : out std_logic_vector(31 downto 0);
    pl_fpd_pll_test_ck_sel_n : in std_logic_vector(2 downto 0);
    pl_fpd_pll_test_fract_clk_sel_n : in std_logic;
    pl_fpd_pll_test_fract_en_n : in std_logic;
    pl_fpd_pll_test_mux_sel : in std_logic_vector(1 downto 0);
    pl_fpd_pll_test_sel : in std_logic_vector(3 downto 0);
    fmio_char_gem_selection : in std_logic_vector(1 downto 0);
    fmio_char_gem_test_select_n : in std_logic;
    fmio_char_gem_test_input : in std_logic;
    fmio_char_gem_test_output : out std_logic;
    test_ddr2pl_dcd_skewout : out std_logic;
    test_pl2ddr_dcd_sample_pulse : in std_logic;
    test_bscan_en_n : in std_logic;
    test_bscan_tdi : in std_logic;
    test_bscan_updatedr : in std_logic;
    test_bscan_shiftdr : in std_logic;
    test_bscan_reset_tap_b : in std_logic;
    test_bscan_misr_jtag_load : in std_logic;
    test_bscan_intest : in std_logic;
    test_bscan_extest : in std_logic;
    test_bscan_clockdr : in std_logic;
    test_bscan_ac_mode : in std_logic;
    test_bscan_ac_test : in std_logic;
    test_bscan_init_memory : in std_logic;
    test_bscan_mode_c : in std_logic;
    test_bscan_tdo : out std_logic;
    i_dbg_l0_txclk : in std_logic;
    i_dbg_l0_rxclk : in std_logic;
    i_dbg_l1_txclk : in std_logic;
    i_dbg_l1_rxclk : in std_logic;
    i_dbg_l2_txclk : in std_logic;
    i_dbg_l2_rxclk : in std_logic;
    i_dbg_l3_txclk : in std_logic;
    i_dbg_l3_rxclk : in std_logic;
    i_afe_rx_symbol_clk_by_2_pl : in std_logic;
    pl_fpd_spare_0_in : in std_logic;
    pl_fpd_spare_1_in : in std_logic;
    pl_fpd_spare_2_in : in std_logic;
    pl_fpd_spare_3_in : in std_logic;
    pl_fpd_spare_4_in : in std_logic;
    fpd_pl_spare_0_out : out std_logic;
    fpd_pl_spare_1_out : out std_logic;
    fpd_pl_spare_2_out : out std_logic;
    fpd_pl_spare_3_out : out std_logic;
    fpd_pl_spare_4_out : out std_logic;
    pl_lpd_spare_0_in : in std_logic;
    pl_lpd_spare_1_in : in std_logic;
    pl_lpd_spare_2_in : in std_logic;
    pl_lpd_spare_3_in : in std_logic;
    pl_lpd_spare_4_in : in std_logic;
    lpd_pl_spare_0_out : out std_logic;
    lpd_pl_spare_1_out : out std_logic;
    lpd_pl_spare_2_out : out std_logic;
    lpd_pl_spare_3_out : out std_logic;
    lpd_pl_spare_4_out : out std_logic;
    o_dbg_l0_phystatus : out std_logic;
    o_dbg_l0_rxdata : out std_logic_vector(19 downto 0);
    o_dbg_l0_rxdatak : out std_logic_vector(1 downto 0);
    o_dbg_l0_rxvalid : out std_logic;
    o_dbg_l0_rxstatus : out std_logic_vector(2 downto 0);
    o_dbg_l0_rxelecidle : out std_logic;
    o_dbg_l0_rstb : out std_logic;
    o_dbg_l0_txdata : out std_logic_vector(19 downto 0);
    o_dbg_l0_txdatak : out std_logic_vector(1 downto 0);
    o_dbg_l0_rate : out std_logic_vector(1 downto 0);
    o_dbg_l0_powerdown : out std_logic_vector(1 downto 0);
    o_dbg_l0_txelecidle : out std_logic;
    o_dbg_l0_txdetrx_lpback : out std_logic;
    o_dbg_l0_rxpolarity : out std_logic;
    o_dbg_l0_tx_sgmii_ewrap : out std_logic;
    o_dbg_l0_rx_sgmii_en_cdet : out std_logic;
    o_dbg_l0_sata_corerxdata : out std_logic_vector(19 downto 0);
    o_dbg_l0_sata_corerxdatavalid : out std_logic_vector(1 downto 0);
    o_dbg_l0_sata_coreready : out std_logic;
    o_dbg_l0_sata_coreclockready : out std_logic;
    o_dbg_l0_sata_corerxsignaldet : out std_logic;
    o_dbg_l0_sata_phyctrltxdata : out std_logic_vector(19 downto 0);
    o_dbg_l0_sata_phyctrltxidle : out std_logic;
    o_dbg_l0_sata_phyctrltxrate : out std_logic_vector(1 downto 0);
    o_dbg_l0_sata_phyctrlrxrate : out std_logic_vector(1 downto 0);
    o_dbg_l0_sata_phyctrltxrst : out std_logic;
    o_dbg_l0_sata_phyctrlrxrst : out std_logic;
    o_dbg_l0_sata_phyctrlreset : out std_logic;
    o_dbg_l0_sata_phyctrlpartial : out std_logic;
    o_dbg_l0_sata_phyctrlslumber : out std_logic;
    o_dbg_l1_phystatus : out std_logic;
    o_dbg_l1_rxdata : out std_logic_vector(19 downto 0);
    o_dbg_l1_rxdatak : out std_logic_vector(1 downto 0);
    o_dbg_l1_rxvalid : out std_logic;
    o_dbg_l1_rxstatus : out std_logic_vector(2 downto 0);
    o_dbg_l1_rxelecidle : out std_logic;
    o_dbg_l1_rstb : out std_logic;
    o_dbg_l1_txdata : out std_logic_vector(19 downto 0);
    o_dbg_l1_txdatak : out std_logic_vector(1 downto 0);
    o_dbg_l1_rate : out std_logic_vector(1 downto 0);
    o_dbg_l1_powerdown : out std_logic_vector(1 downto 0);
    o_dbg_l1_txelecidle : out std_logic;
    o_dbg_l1_txdetrx_lpback : out std_logic;
    o_dbg_l1_rxpolarity : out std_logic;
    o_dbg_l1_tx_sgmii_ewrap : out std_logic;
    o_dbg_l1_rx_sgmii_en_cdet : out std_logic;
    o_dbg_l1_sata_corerxdata : out std_logic_vector(19 downto 0);
    o_dbg_l1_sata_corerxdatavalid : out std_logic_vector(1 downto 0);
    o_dbg_l1_sata_coreready : out std_logic;
    o_dbg_l1_sata_coreclockready : out std_logic;
    o_dbg_l1_sata_corerxsignaldet : out std_logic;
    o_dbg_l1_sata_phyctrltxdata : out std_logic_vector(19 downto 0);
    o_dbg_l1_sata_phyctrltxidle : out std_logic;
    o_dbg_l1_sata_phyctrltxrate : out std_logic_vector(1 downto 0);
    o_dbg_l1_sata_phyctrlrxrate : out std_logic_vector(1 downto 0);
    o_dbg_l1_sata_phyctrltxrst : out std_logic;
    o_dbg_l1_sata_phyctrlrxrst : out std_logic;
    o_dbg_l1_sata_phyctrlreset : out std_logic;
    o_dbg_l1_sata_phyctrlpartial : out std_logic;
    o_dbg_l1_sata_phyctrlslumber : out std_logic;
    o_dbg_l2_phystatus : out std_logic;
    o_dbg_l2_rxdata : out std_logic_vector(19 downto 0);
    o_dbg_l2_rxdatak : out std_logic_vector(1 downto 0);
    o_dbg_l2_rxvalid : out std_logic;
    o_dbg_l2_rxstatus : out std_logic_vector(2 downto 0);
    o_dbg_l2_rxelecidle : out std_logic;
    o_dbg_l2_rstb : out std_logic;
    o_dbg_l2_txdata : out std_logic_vector(19 downto 0);
    o_dbg_l2_txdatak : out std_logic_vector(1 downto 0);
    o_dbg_l2_rate : out std_logic_vector(1 downto 0);
    o_dbg_l2_powerdown : out std_logic_vector(1 downto 0);
    o_dbg_l2_txelecidle : out std_logic;
    o_dbg_l2_txdetrx_lpback : out std_logic;
    o_dbg_l2_rxpolarity : out std_logic;
    o_dbg_l2_tx_sgmii_ewrap : out std_logic;
    o_dbg_l2_rx_sgmii_en_cdet : out std_logic;
    o_dbg_l2_sata_corerxdata : out std_logic_vector(19 downto 0);
    o_dbg_l2_sata_corerxdatavalid : out std_logic_vector(1 downto 0);
    o_dbg_l2_sata_coreready : out std_logic;
    o_dbg_l2_sata_coreclockready : out std_logic;
    o_dbg_l2_sata_corerxsignaldet : out std_logic;
    o_dbg_l2_sata_phyctrltxdata : out std_logic_vector(19 downto 0);
    o_dbg_l2_sata_phyctrltxidle : out std_logic;
    o_dbg_l2_sata_phyctrltxrate : out std_logic_vector(1 downto 0);
    o_dbg_l2_sata_phyctrlrxrate : out std_logic_vector(1 downto 0);
    o_dbg_l2_sata_phyctrltxrst : out std_logic;
    o_dbg_l2_sata_phyctrlrxrst : out std_logic;
    o_dbg_l2_sata_phyctrlreset : out std_logic;
    o_dbg_l2_sata_phyctrlpartial : out std_logic;
    o_dbg_l2_sata_phyctrlslumber : out std_logic;
    o_dbg_l3_phystatus : out std_logic;
    o_dbg_l3_rxdata : out std_logic_vector(19 downto 0);
    o_dbg_l3_rxdatak : out std_logic_vector(1 downto 0);
    o_dbg_l3_rxvalid : out std_logic;
    o_dbg_l3_rxstatus : out std_logic_vector(2 downto 0);
    o_dbg_l3_rxelecidle : out std_logic;
    o_dbg_l3_rstb : out std_logic;
    o_dbg_l3_txdata : out std_logic_vector(19 downto 0);
    o_dbg_l3_txdatak : out std_logic_vector(1 downto 0);
    o_dbg_l3_rate : out std_logic_vector(1 downto 0);
    o_dbg_l3_powerdown : out std_logic_vector(1 downto 0);
    o_dbg_l3_txelecidle : out std_logic;
    o_dbg_l3_txdetrx_lpback : out std_logic;
    o_dbg_l3_rxpolarity : out std_logic;
    o_dbg_l3_tx_sgmii_ewrap : out std_logic;
    o_dbg_l3_rx_sgmii_en_cdet : out std_logic;
    o_dbg_l3_sata_corerxdata : out std_logic_vector(19 downto 0);
    o_dbg_l3_sata_corerxdatavalid : out std_logic_vector(1 downto 0);
    o_dbg_l3_sata_coreready : out std_logic;
    o_dbg_l3_sata_coreclockready : out std_logic;
    o_dbg_l3_sata_corerxsignaldet : out std_logic;
    o_dbg_l3_sata_phyctrltxdata : out std_logic_vector(19 downto 0);
    o_dbg_l3_sata_phyctrltxidle : out std_logic;
    o_dbg_l3_sata_phyctrltxrate : out std_logic_vector(1 downto 0);
    o_dbg_l3_sata_phyctrlrxrate : out std_logic_vector(1 downto 0);
    o_dbg_l3_sata_phyctrltxrst : out std_logic;
    o_dbg_l3_sata_phyctrlrxrst : out std_logic;
    o_dbg_l3_sata_phyctrlreset : out std_logic;
    o_dbg_l3_sata_phyctrlpartial : out std_logic;
    o_dbg_l3_sata_phyctrlslumber : out std_logic;
    dbg_path_fifo_bypass : out std_logic;
    i_afe_pll_pd_hs_clock_r : in std_logic;
    i_afe_mode : in std_logic;
    i_bgcal_afe_mode : in std_logic;
    o_afe_cmn_calib_comp_out : out std_logic;
    i_afe_cmn_bg_enable_low_leakage : in std_logic;
    i_afe_cmn_bg_iso_ctrl_bar : in std_logic;
    i_afe_cmn_bg_pd : in std_logic;
    i_afe_cmn_bg_pd_bg_ok : in std_logic;
    i_afe_cmn_bg_pd_ptat : in std_logic;
    i_afe_cmn_calib_en_iconst : in std_logic;
    i_afe_cmn_calib_enable_low_leakage : in std_logic;
    i_afe_cmn_calib_iso_ctrl_bar : in std_logic;
    o_afe_pll_dco_count : out std_logic_vector(12 downto 0);
    o_afe_pll_clk_sym_hs : out std_logic;
    o_afe_pll_fbclk_frac : out std_logic;
    o_afe_rx_pipe_lfpsbcn_rxelecidle : out std_logic;
    o_afe_rx_pipe_sigdet : out std_logic;
    o_afe_rx_symbol : out std_logic_vector(19 downto 0);
    o_afe_rx_symbol_clk_by_2 : out std_logic;
    o_afe_rx_uphy_save_calcode : out std_logic;
    o_afe_rx_uphy_startloop_buf : out std_logic;
    o_afe_rx_uphy_rx_calib_done : out std_logic;
    i_afe_rx_rxpma_rstb : in std_logic;
    i_afe_rx_uphy_restore_calcode_data : in std_logic_vector(7 downto 0);
    i_afe_rx_pipe_rxeqtraining : in std_logic;
    i_afe_rx_iso_hsrx_ctrl_bar : in std_logic;
    i_afe_rx_iso_lfps_ctrl_bar : in std_logic;
    i_afe_rx_iso_sigdet_ctrl_bar : in std_logic;
    i_afe_rx_hsrx_clock_stop_req : in std_logic;
    o_afe_rx_uphy_save_calcode_data : out std_logic_vector(7 downto 0);
    o_afe_rx_hsrx_clock_stop_ack : out std_logic;
    o_afe_pg_avddcr : out std_logic;
    o_afe_pg_avddio : out std_logic;
    o_afe_pg_dvddcr : out std_logic;
    o_afe_pg_static_avddcr : out std_logic;
    o_afe_pg_static_avddio : out std_logic;
    i_pll_afe_mode : in std_logic;
    i_afe_pll_coarse_code : in std_logic_vector(10 downto 0);
    i_afe_pll_en_clock_hs_div2 : in std_logic;
    i_afe_pll_fbdiv : in std_logic_vector(15 downto 0);
    i_afe_pll_load_fbdiv : in std_logic;
    i_afe_pll_pd : in std_logic;
    i_afe_pll_pd_pfd : in std_logic;
    i_afe_pll_rst_fdbk_div : in std_logic;
    i_afe_pll_startloop : in std_logic;
    i_afe_pll_v2i_code : in std_logic_vector(5 downto 0);
    i_afe_pll_v2i_prog : in std_logic_vector(4 downto 0);
    i_afe_pll_vco_cnt_window : in std_logic;
    i_afe_rx_mphy_gate_symbol_clk : in std_logic;
    i_afe_rx_mphy_mux_hsb_ls : in std_logic;
    i_afe_rx_pipe_rx_term_enable : in std_logic;
    i_afe_rx_uphy_biasgen_iconst_core_mirror_enable : in std_logic;
    i_afe_rx_uphy_biasgen_iconst_io_mirror_enable : in std_logic;
    i_afe_rx_uphy_biasgen_irconst_core_mirror_enable : in std_logic;
    i_afe_rx_uphy_enable_cdr : in std_logic;
    i_afe_rx_uphy_enable_low_leakage : in std_logic;
    i_afe_rx_rxpma_refclk_dig : in std_logic;
    i_afe_rx_uphy_hsrx_rstb : in std_logic;
    i_afe_rx_uphy_pdn_hs_des : in std_logic;
    i_afe_rx_uphy_pd_samp_c2c : in std_logic;
    i_afe_rx_uphy_pd_samp_c2c_eclk : in std_logic;
    i_afe_rx_uphy_pso_clk_lane : in std_logic;
    i_afe_rx_uphy_pso_eq : in std_logic;
    i_afe_rx_uphy_pso_hsrxdig : in std_logic;
    i_afe_rx_uphy_pso_iqpi : in std_logic;
    i_afe_rx_uphy_pso_lfpsbcn : in std_logic;
    i_afe_rx_uphy_pso_samp_flops : in std_logic;
    i_afe_rx_uphy_pso_sigdet : in std_logic;
    i_afe_rx_uphy_restore_calcode : in std_logic;
    i_afe_rx_uphy_run_calib : in std_logic;
    i_afe_rx_uphy_rx_lane_polarity_swap : in std_logic;
    i_afe_rx_uphy_startloop_pll : in std_logic;
    i_afe_rx_uphy_hsclk_division_factor : in std_logic_vector(1 downto 0);
    i_afe_rx_uphy_rx_pma_opmode : in std_logic_vector(7 downto 0);
    i_afe_tx_enable_hsclk_division : in std_logic_vector(1 downto 0);
    i_afe_tx_enable_ldo : in std_logic;
    i_afe_tx_enable_ref : in std_logic;
    i_afe_tx_enable_supply_hsclk : in std_logic;
    i_afe_tx_enable_supply_pipe : in std_logic;
    i_afe_tx_enable_supply_serializer : in std_logic;
    i_afe_tx_enable_supply_uphy : in std_logic;
    i_afe_tx_hs_ser_rstb : in std_logic;
    i_afe_tx_hs_symbol : in std_logic_vector(19 downto 0);
    i_afe_tx_mphy_tx_ls_data : in std_logic;
    i_afe_tx_pipe_tx_enable_idle_mode : in std_logic_vector(1 downto 0);
    i_afe_tx_pipe_tx_enable_lfps : in std_logic_vector(1 downto 0);
    i_afe_tx_pipe_tx_enable_rxdet : in std_logic;
    i_afe_TX_uphy_txpma_opmode : in std_logic_vector(7 downto 0);
    i_afe_TX_pmadig_digital_reset_n : in std_logic;
    i_afe_TX_serializer_rst_rel : in std_logic;
    i_afe_TX_pll_symb_clk_2 : in std_logic;
    i_afe_TX_ana_if_rate : in std_logic_vector(1 downto 0);
    i_afe_TX_en_dig_sublp_mode : in std_logic;
    i_afe_TX_LPBK_SEL : in std_logic_vector(2 downto 0);
    i_afe_TX_iso_ctrl_bar : in std_logic;
    i_afe_TX_ser_iso_ctrl_bar : in std_logic;
    i_afe_TX_lfps_clk : in std_logic;
    i_afe_TX_serializer_rstb : in std_logic;
    o_afe_TX_dig_reset_rel_ack : out std_logic;
    o_afe_TX_pipe_TX_dn_rxdet : out std_logic;
    o_afe_TX_pipe_TX_dp_rxdet : out std_logic;
    i_afe_tx_pipe_tx_fast_est_common_mode : in std_logic;
    o_dbg_l0_txclk : out std_logic;
    o_dbg_l0_rxclk : out std_logic;
    o_dbg_l1_txclk : out std_logic;
    o_dbg_l1_rxclk : out std_logic;
    o_dbg_l2_txclk : out std_logic;
    o_dbg_l2_rxclk : out std_logic;
    o_dbg_l3_txclk : out std_logic;
    o_dbg_l3_rxclk : out std_logic
  );
end component;

component zynq_ultra_ps_e is
  port(
    ps_in        : in    pl2ps_t;
    ps_out       : out   ps2pl_t;
    m_axi_hp_in  : in    m_axi_hp_in_array_t(0 to C_M_AXI_HP_COUNT-1);
    m_axi_hp_out : out   m_axi_hp_out_array_t(0 to C_M_AXI_HP_COUNT-1);
    s_axi_hp_in  : in    s_axi_hp_in_array_t(0 to C_S_AXI_HP_COUNT-1);
    s_axi_hp_out : out   s_axi_hp_out_array_t(0 to C_S_AXI_HP_COUNT-1)
    );
end component zynq_ultra_ps_e;
end package zynq_ultra_pkg;
