../../../bias_param.rcc/target-2-linux-c6-x86_64/generics.vhd