-- The SDP Sender, to take data from a WSI port, and put it in memory, making it available
-- for someone to read it out and acknowledge that reading.

library IEEE, ocpi, util, bsv, sdp;
use IEEE.std_logic_1164.all, ieee.numeric_std.all, ocpi.types.all, ocpi.util.all, sdp.all;
architecture rtl of sdp_send_worker is
  -- Local worker constants
  constant sdp_width_c    : natural := to_integer(sdp_width);
  constant memory_depth_c : natural := to_integer(memory_bytes) / (sdp_width_c * 4);
  constant addr_width_c   : natural := width_for_max(memory_depth_c - 1);
  constant max_buffers_c  : natural := to_integer(max_buffers);
  constant addr_shift_c   : natural := width_for_max(sdp_width_c * 4 - 1);
  constant count_width_c  : natural := width_for_max(max_buffers_c);
  constant nbytes_width_c : natural := width_for_max(sdp_width_c * 4); -- nbytes in frame
  constant max_remotes_c  : natural := to_integer(max_remotes);

  -- Metadata (internal) FIFO definitions
  constant meta_length_c  : natural := 0;
  constant meta_length_width_c : natural := 23;
  constant meta_eof_c     : natural := meta_length_c + meta_length_width_c;
  constant meta_opcode_c  : natural := meta_eof_c + 1;
  constant meta_opcode_width_c  : natural := 8;
  type metadata_t is record
    length : unsigned(meta_length_width_c-1 downto 0); -- bytes
    eof    : bool_t;
    opcode : std_logic_vector(meta_opcode_width_c-1 downto 0);
  end record metadata_t;
  constant metawidth_c : integer := meta_length_width_c + 1 + meta_opcode_width_c;
  constant meta_ndws_c : integer := (metawidth_c + dword_size - 1) / dword_size;
  function meta2slv(meta : metadata_t) return std_logic_vector is
  begin
    return meta.opcode & slv(meta.eof) & slv(meta.length);
  end meta2slv;
  function slv2meta(s : std_logic_vector(metawidth_c-1 downto 0)) return metadata_t is
    variable m : metadata_t;
  begin
    m.length := unsigned(s(meta_length_width_c-1 downto 0));
    m.eof    := s(meta_length_c);
    m.opcode := s(s'left downto meta_eof_c + 1);
    return m;
  end slv2meta;

  subtype remote_idx_t is unsigned(width_for_max(max_remotes_c - 1) - 1 downto 0);

  -- Flag/doorbell Sync FIFO definitions
  signal flag_enq       : bool_t;
  signal flag_in_remote : remote_idx_t;
  signal flag_not_full  : std_logic;
  signal flag_deq       : bool_t;
  signal flag_out_slv   : std_logic_vector(remote_idx_t'range);
  signal flag_out       : natural;
  signal flag_not_empty : std_logic;

  -- Metadata definitions for the SDP side
  constant sdp_meta_ndws_c : natural := 2;

  -- Convenience data types
  subtype buffer_count_t is unsigned(count_width_c - 1 downto 0);
  subtype bram_addr_t is unsigned(addr_width_c-1 downto 0);

  -- Definitions for remote accesses
  constant sdp_whole_addr_bits_c : integer := sdp.sdp.addr_width + sdp.sdp.node_width;
  subtype sdp_whole_addr_t is unsigned(sdp_whole_addr_bits_c-1 downto 0);
  -- Dynamic state of a remote destination (static state is in properties)
  type remote_t is record
    index     : buffer_count_t; -- which remote buffer are we sending to?
    empty     : buffer_count_t; -- how many remote buffers are empty?
    data_addr : sdp_whole_addr_t;
    meta_addr : sdp_whole_addr_t;
    flag_addr : sdp_whole_addr_t;
  end record remote_t;
  type remote_array_t is array(0 to max_remotes_c-1) of remote_t;
  signal sdp_remotes : remote_array_t;

  -- Combinatorial signals
  signal can_take          : bool_t;
  signal will_write        : bool_t;
  signal max_offset        : bram_addr_t;
  signal next_buffer_addr  : bram_addr_t;
  signal bram_addr         : bram_addr_t;
  signal bram_addr_actual  : bram_addr_t;
  signal bad_write         : bool_t;
  signal nbytes            : unsigned(nbytes_width_c-1 downto 0);
  -- Registered signals
  ---- WSI buffer filling pointers
  signal buffer_offset_r   : bram_addr_t;    -- offset in current buffer
  signal buffer_index_r    : buffer_count_t;
  signal buffer_addr_r     : bram_addr_t;    -- base of current buffer
  signal buffer_avail_r    : buffer_count_t; -- how local many buffers are empty?
  signal buffer_consumed   : bool_t;         -- pulse for buffer consumption from sdp side
  ---- Metadata management
  signal md_r              : ulong_array_t(0 to max_Buffers_c - 1); -- readback property
  signal md_in             : metadata_t;
  signal md_out            : metadata_t;
  signal md_out_slv        : std_logic_vector(metawidth_c-1 downto 0);
  signal md_enq            : bool_t;
  signal md_deq            : std_logic;
  signal md_not_empty      : std_logic;
  signal md_not_full       : std_logic;
  -- ndws is rounded up so needs ONE fewer bits, not TWO
  signal md_out_ndws       : unsigned(meta_length_width_c-2 downto 0);

  -- SDP back side --
  signal bramb_addr             : bram_addr_t;
  signal bramb_addr_r           : bram_addr_t;
  signal bramb_out              : std_logic_vector(sdp_width_c*32-1 downto 0);
  signal sdp_out_r              : std_logic_vector(sdp_width_c*32-1 downto 0);
  signal sdp_out_valid_r        : bool_t;
  signal sdp_segment_count_r    : sdp.sdp.count_t;
  signal sdp_last_in_segment    : bool_t;
  -- State that changes for each msg
  signal sdp_msg_idx_r          : buffer_count_t;
  signal sdp_next_msg_addr      : bram_addr_t;
  signal sdp_msg_addr_r         : bram_addr_t;
  -- State that changes for each remote
  type sdp_phase_t is (idle_e, data_e, meta_e, flag_e, between_remotes_e);
  signal sdp_remote_phase_r     : sdp_phase_t;
  subtype meta_dw_count_t is unsigned(meta_length_width_c-2 downto 0);
  signal sdp_msg_dws_left_r     : meta_dw_count_t;
  signal sdp_remote_idx_r       : remote_idx_t;
  signal sdp_last_remote        : remote_idx_t;
  -- State that changed for each segment
  signal sdp_segment_addr_r     : sdp_whole_addr_t;
  signal sdp_whole_addr         : sdp_whole_addr_t;
  signal sdp_segment_dws_left_r : meta_dw_count_t;

  ---- Global state
  signal overflow_r        : bool_t; -- tried to write past the end of the buffer
  signal operating_r       : bool_t; -- were we operating in the last cycle?
  signal ctl_reset_n       : std_logic;
  signal sdp_reset_n       : std_logic;
  function be2bytes (be    : std_logic_vector) return unsigned is
  begin
    for i in 0 to be'length-1 loop
      if be(i) = '0' then
        return to_unsigned(i, nbytes_width_c);
      end if;
    end loop;
    return to_unsigned(be'length, nbytes_width_c);
  end be2bytes;
begin
  ctl_reset_n        <= not ctl_in.reset;
  bram_addr          <= buffer_addr_r + buffer_offset_r;
  bram_addr_actual   <= bram_addr(addr_width_c-1 downto 0);
  next_buffer_addr   <= buffer_addr_r +
                        props_in.buffer_size(bram_addr_t'left + addr_shift_c
                                             downto addr_shift_c);
  can_take           <= to_bool(operating_r and not its(overflow_r) and md_not_full and buffer_avail_r /= 0);
  will_write         <= can_take and in_in.ready and in_in.valid and not bad_write;
  max_offset         <= props_in.buffer_size(bram_addr_t'left + 2 downto 2) - 1;
  bad_write          <= to_bool((buffer_offset_r > max_offset) or
                                (bram_addr >= memory_depth_c - 1));
  in_out.take        <= can_take and in_in.ready and
                        (will_write or md_enq or (in_in.som and not in_in.valid));
  ctl_out.finished   <= overflow_r;
  props_out.overflow <= overflow_r;
  props_out.sdp_id   <= resize(sdp_in.id, props_out.sdp_id'length);
  props_out.raw.done <= btrue;
  nbytes <= be2bytes(in_in.byte_enable) when its(in_in.valid) else (others => '0');
  md_in.length <= (resize(buffer_offset_r, meta_length_width_c) sll addr_shift_c) + nbytes;
  md_in.eof    <= not in_in.eom and not in_in.som and not in_in.valid;
  md_in.opcode <= in_in.opcode;
  md_enq <= to_bool(its(can_take) and in_in.ready and in_in.eom and
                          its((not in_in.valid) or not bad_write));
  -- Instance the message data BRAM
  -- Since the BRAM is single cycle, there is no handshake.
  bram : component util.util.BRAM2
    generic map(PIPELINED  => 0,
                ADDR_WIDTH => addr_width_c,
                DATA_WIDTH => sdp_width_c * 32,
                MEMSIZE    => memory_depth_c)
    port map   (CLKA       => ctl_in.clk,
                ENA        => '1',
                WEA        => will_write,
                ADDRA      => std_logic_vector(bram_addr_actual),
                DIA        => in_in.data,
                DOA        => open,
                CLKB       => sdp_in.clk,
                ENB        => '1',
                WEB        => '0',
                ADDRB      => std_logic_vector(bramb_addr),
                DIB        => slv0(sdp_width_c*32),
                DOB        => bramb_out);
  
  metafifo : component bsv.bsv.SyncFIFO
   generic map(dataWidth    => metawidth_c,
               depth        => roundup_2_power_of_2(max_buffers_c), -- must be power of 2
               indxWidth    => width_for_max(roundup_2_power_of_2(max_buffers_c)-1))
   port map   (sCLK         => ctl_in.clk,
               sRST         => ctl_reset_n,
               dCLK         => sdp_in.clk,
               sENQ         => std_logic(md_enq),
               sD_IN        => meta2slv(md_in),
               sFULL_N      => md_not_full,
               dDEQ         => md_deq,
               dD_OUT       => md_out_slv,
               dEMPTY_N     => md_not_empty);

  -- A sync fifo to carry doorbells to the SDP clock domain
  flagfifo : component bsv.bsv.SyncFIFO
   generic map(dataWidth    => remote_idx_t'length,
               depth        => 2, -- must be power of 2
               indxWidth    => width_for_max(2-1))
   port map   (sCLK         => ctl_in.clk, -- maybe syncfifo later
               sRST         => ctl_reset_n,
               dCLK         => sdp_in.clk,
               sENQ         => std_logic(flag_enq),
               sD_IN        => std_logic_vector(flag_in_remote),
               sFULL_N      => flag_not_full,
               dDEQ         => flag_deq,
               dD_OUT       => flag_out_slv,
               dEMPTY_N     => flag_not_empty);

  -- A sync pulse to carry buffer consumption events
  cpulse: component bsv.bsv.SyncPulse
    port map  (sCLK         => sdp_in.clk,
               sRST         => sdp_reset_n,
               dCLK         => ctl_in.clk,
               sEN          => md_deq,
               dPulse       => buffer_consumed);
  -- source side
  flag_enq       <= props_in.raw.is_write; -- the only raw thing written
  flag_in_remote <= props_in.raw.address(flag_in_remote'length-1+2 downto 2); -- ulongs/dws
  -- destination side
  flag_out       <= to_integer(remote_idx_t(flag_out_slv));
  flag_deq       <= flag_not_empty; -- output of FIFO always processed immediately

  -- the process going from wsi into the data bram and metadata fifo
  wsi2bram : process(ctl_in.clk)
  begin
    if rising_edge(ctl_in.clk) then
      if ctl_in.reset = '1' then
        buffer_offset_r <= (others => '0');
        buffer_index_r  <= (others => '0');
        buffer_addr_r   <= (others => '0');
        operating_r     <= bfalse;
        overflow_r      <= bfalse;
      elsif not operating_r then
        -- initialization on first transition to operating.  poor man's "start".
        if its(ctl_in.is_operating) then
          operating_r   <= btrue;
          if props_in.buffer_size > memory_bytes then
            overflow_r <= btrue;
          end if;
        end if;
        buffer_avail_r <= resize(props_in.buffer_count, buffer_avail_r'length);
      elsif not ctl_in.is_operating then
        operating_r <= bfalse;
      else
        if md_enq and not its(buffer_consumed) then
          buffer_avail_r <= buffer_avail_r - 1;
        end if;
        if buffer_consumed and not its(md_enq) then
          buffer_avail_r <= buffer_avail_r + 1;
        end if;
        if props_in.raw.is_write and not flag_not_full = '1' then
          overflow_r <= btrue; -- this is really a debug thing.  Should not happen.
        end if;
        if can_take and in_in.ready then
          if its(in_in.valid) then
            if its(bad_write) then
              overflow_r <= btrue; -- this should be sticky
            end if;
            buffer_offset_r <= buffer_offset_r + 1;
          end if;
          if in_in.eom or its(not in_in.eom and not in_in.som and not in_in.valid) then
            buffer_offset_r   <= (others => '0');
            if buffer_index_r = props_in.buffer_count - 1 then
              buffer_index_r  <= (others => '0');
              buffer_addr_r   <= (others => '0');
            else
              buffer_index_r  <= buffer_index_r + 1;
              buffer_addr_r   <= next_buffer_addr;
            end if;
          end if; -- eom
        end if; -- cantake and ready
      end if; -- operating
    end if; -- rising edge
  end process;

  --------------------------------------------------------------------------------
  -- BRAM to SDP signals and process, in the clock domain from the SDP.
  sdp_reset_n         <= not sdp_in.reset;
  sdp_last_remote     <= resize(props_in.remote_count -1, remote_idx_t'length);
  md_out              <= slv2meta(md_out_slv);
  md_out_ndws         <= resize((md_out.length + dword_bytes - 1) srl 2, md_out_ndws'length);
  md_deq              <= operating_r and md_not_empty and sdp_in.sdp.ready and
                         to_bool(sdp_remote_phase_r = flag_e) and
                         to_bool(sdp_remote_idx_r = sdp_last_remote);
  sdp_last_in_segment <= to_bool(sdp_segment_dws_left_r = 0);
  -- What is the address of the next message in BRAM
  sdp_next_msg_addr   <= sdp_msg_addr_r  when sdp_remote_idx_r /= sdp_last_remote else
                         (others => '0') when sdp_msg_idx_r = props_in.buffer_count - 1 else
                         sdp_msg_addr_r + props_in.buffer_size(bram_addr_t'left + addr_shift_c
                                                               downto addr_shift_c);
  -- The BRAM address must be pipelined (early).
  bramb_addr          <= sdp_next_msg_addr when sdp_remote_phase_r /= data_e else
                         sdp_msg_addr_r when its(sdp_last_in_segment) else
                         bramb_addr_r;
  -- Drive SDP outputs
  sdp_out.sdp.header.op    <= sdp.sdp.write_e;          -- we are only writing
  sdp_out.sdp.header.xid   <= (others => '0');  -- since we are writing, no xid necessary
  sdp_out.sdp.header.lead  <= (others => '0');  -- we are always aligned on a DW
  sdp_out.sdp.header.trail <= (others => '0');  -- we always send whole DWs
  sdp_out.sdp.header.count <= sdp_segment_count_r;
  with sdp_remote_phase_r select sdp_whole_addr <=
    sdp_segment_addr_r                                  when data_e,
    sdp_remotes(to_integer(sdp_remote_idx_r)).meta_addr when meta_e,
    sdp_remotes(to_integer(sdp_remote_idx_r)).flag_addr when flag_e | idle_e | between_remotes_e;
  sdp_out.sdp.header.node  <= sdp_whole_addr(sdp_whole_addr_bits_c-1 downto sdp.sdp.addr_width);
  sdp_out.sdp.header.addr  <= sdp_whole_addr(sdp.sdp.addr_width-1 downto 0);
  sdp_out.sdp.eom          <= sdp_last_in_segment;
  sdp_out.sdp.valid        <= to_bool(sdp_remote_phase_r /= idle_e);
  sdp_out.sdp.ready        <= bfalse;     -- we are write-only, never accepting an inbound frame
g0: for i in 0 to sdp_width_c-1 generate
    sdp_out_data(i) <= sdp_out_r((i+1)*dword_size-1 downto i*dword_size)
                       when its(sdp_out_valid_r) else
                       bramb_out((i+1)*dword_size-1 downto i*dword_size);
  end generate g0;

  -- The process that takes messages from BRAM and pushes them to the SDP,
  ---- trying to avoid any dead cycles except one at the start of the message
  ---- sending data(except for ZLM), metadata, flag transfers
  ---- breaking up the data messages into SDP-required segments
  bram2sdp : process(sdp_in.clk)
    variable r : natural;
    variable started_remote : boolean;
    impure function remote_is_ready(r : natural) return boolean is
    begin
      return sdp_remotes(r).empty /= 0 or (flag_not_empty = '1' and flag_out = r);
    end remote_is_ready;
    procedure begin_segment(ndws_left : meta_dw_count_t) is
      variable ndws : unsigned(ndws_left'range);
    begin
      if ndws_left > sdp.sdp.max_segment_dws then
        ndws :=  to_unsigned(sdp.sdp.max_segment_dws, ndws'length);
      else
        ndws :=  ndws_left;
      end if;
      if ndws <= sdp_width then
        sdp_segment_dws_left_r <= (others => '0');
      else
        sdp_segment_dws_left_r <= ndws - sdp_width;
      end if;
      sdp_msg_dws_left_r     <= ndws_left - ndws; -- this does no harm in non-data phases
      sdp_segment_count_r    <= resize(ndws - 1, sdp_segment_count_r'length);
    end procedure begin_segment;
    -- Start a segment, given how many DWs are left in the message,
    -- and set the left-in-segment, left-in-message, and segment header count
    procedure begin_meta is
      variable meta :std_logic_vector(39 downto 0)
        := md_out.opcode & std_logic_vector(resize(md_out.length, 32));
    begin
      sdp_out_r <= std_logic_vector(meta(sdp_out_r'range));
      sdp_remote_phase_r <= meta_e;
      sdp_out_valid_r    <= btrue;
      begin_segment(to_unsigned(sdp_meta_ndws_c, meta_dw_count_t'length));
    end procedure begin_meta;
    -- initialization for sending the current message to the indicated remote
    procedure begin_remote is
      variable data_addr : sdp_whole_addr_t;
      variable meta_addr : sdp_whole_addr_t;
      variable flag_addr : sdp_whole_addr_t;
    begin
      started_remote := true;
      sdp_remote_idx_r   <= to_unsigned(r, sdp_remote_idx_r'length);
      if sdp_remotes(r).index = 0 then
        data_addr := props_in.remote_data_addr(r)(data_addr'left+2 downto 2);
        meta_addr := props_in.remote_meta_addr(r)(meta_addr'left+2 downto 2);
        flag_addr := props_in.remote_flag_addr(r)(flag_addr'left+2 downto 2);
      else
        data_addr := sdp_remotes(r).data_addr +
                     resize(props_in.remote_data_pitch(r)(ulong_t'left downto 2),
                            sdp_whole_addr_t'length);
        meta_addr := sdp_remotes(r).meta_addr +
                     resize(props_in.remote_meta_pitch(r)(ulong_t'left downto 2),
                            sdp_whole_addr_t'length);
        flag_addr := sdp_remotes(r).flag_addr +
                     resize(props_in.remote_flag_pitch(r)(ulong_t'left downto 2),
                            sdp_whole_addr_t'length);
      end if;
      sdp_remotes(r).data_addr <= data_addr;
      sdp_remotes(r).meta_addr <= meta_addr;
      sdp_remotes(r).flag_addr <= flag_addr;
      if sdp_remotes(r).index = props_in.remote_buffer_count(r) - 1 then
        sdp_remotes(r).index <= (others => '0');
      else
        sdp_remotes(r).index <= sdp_remotes(r).index + 1;
      end if;
      if md_out_ndws = 0 then
        begin_meta;
        sdp_segment_addr_r <= meta_addr;
      else
        sdp_remote_phase_r <= data_e;
        sdp_segment_addr_r <= data_addr;
        sdp_out_r          <= bramb_out;
        sdp_out_valid_r    <= btrue;
        begin_segment(md_out_ndws);
      end if;
    end procedure begin_remote;
  begin
    r              := to_integer(sdp_remote_idx_r);
    started_remote := false;
    if rising_edge(sdp_in.clk) then
      if its(sdp_in.reset) then
        -- Reset state for remotes
        for r in 0 to max_remotes_c - 1 loop
          sdp_remotes(r).index <= (others => '0');
        end loop;
        sdp_remote_phase_r <= idle_e;
        sdp_remote_idx_r   <= (others => '0');
      elsif not operating_r then
        -- reset state that depends on properties
        for r in 0 to max_remotes_c - 1 loop
          sdp_remotes(r).empty <= resize(props_in.remote_buffer_count(r),buffer_count_t'length);
        end loop;
        sdp_msg_idx_r <= resize(props_in.buffer_count - 1, sdp_msg_idx_r'length);
      else
        if md_not_empty = '1' then
          if sdp_remote_phase_r = idle_e then
            if remote_is_ready(0) then
              -- We are starting to send a message to all remotes.  bram addr was already valid
              sdp_msg_addr_r <= sdp_next_msg_addr;
              bramb_addr_r   <= sdp_next_msg_addr + 1;
              begin_remote;
            end if;
          elsif sdp_remote_phase_r = between_remotes_e then
            if remote_is_ready(r) then
              begin_remote;
            end if;
          elsif its(sdp_in.sdp.ready) then
            if sdp_segment_dws_left_r /= 0 then
              -- continue the segment
              case sdp_remote_phase_r is
                when data_e =>
                  bramb_addr_r <= bramb_addr + 1; -- this is irrelevant to meta and flag phases
                  sdp_out_valid_r <= bfalse;
                when meta_e => -- must be single word width
                  sdp_out_r <= std_logic_vector(resize(unsigned(md_out.opcode), sdp_out_r'length));
                  sdp_out_valid_r <= btrue;
                when others => null;
              end case;
              sdp_segment_dws_left_r <= sdp_segment_dws_left_r - sdp_width_c;
            else
              -- end the segment
              case sdp_remote_phase_r is
                when data_e =>
                  if sdp_msg_dws_left_r /= 0 then
                    begin_segment(sdp_msg_dws_left_r);
                  else
                    begin_meta;
                  end if;
                when meta_e =>
                  sdp_segment_count_r <= (others => '0');
                  sdp_remote_phase_r  <= flag_e;
                  sdp_out_r           <= std_logic_vector(to_unsigned(1, sdp_out_r'length));
                  -- Advance the buffer pointer here (not in flag_e) to pipeline the bram address
                  if r = sdp_last_remote then
                    if sdp_msg_idx_r = props_in.buffer_count - 1 then
                      sdp_msg_idx_r    <= (others => '0');
                    else
                      sdp_msg_idx_r    <= sdp_msg_idx_r + 1;
                    end if;
                  end if;
                when flag_e =>
                  -- end of transferring a message to a remote
                  if r = sdp_last_remote then
                    sdp_remote_phase_r <= idle_e; -- our one idle cycle per message
                    sdp_remote_idx_r   <= (others => '0');
                  else
                    -- move on to the next remote with the same message
                    r := r + 1;
                    bramb_addr_r <= sdp_msg_addr_r + 1;
                    if remote_is_ready(r) then
                      begin_remote;
                    else
                      sdp_remote_idx_r   <= to_unsigned(r, sdp_remote_idx_r'length);
                      sdp_remote_phase_r <= between_remotes_e;
                    end if;
                  end if;
                when others => null;
              end case;
            end if; -- if/else end of segment
          end if; -- if/else idle
        end if; -- message available in fifo 
        -- Process doorbells
        if flag_not_empty = '1' and not (started_remote and flag_out = r) then
          sdp_remotes(flag_out).empty <= sdp_remotes(flag_out).empty + 1;
        end if;
        if started_remote and not (flag_not_empty = '1' and flag_out = r) then
          sdp_remotes(r).empty <= sdp_remotes(r).empty - 1;
        end if;
      end if; -- if/else reset/operating
    end if; -- if rising edge
  end process;
end architecture rtl;
