-- THIS FILE WAS ORIGINALLY GENERATED ON Tue Apr 16 15:05:54 2013 EDT
-- BASED ON THE FILE: bias_vhdl1.xml
-- YOU *ARE* EXPECTED TO EDIT IT
-- This file initially contains the architecture skeleton for worker: bias_vhdl1

library IEEE; use IEEE.std_logic_1164.all; use ieee.numeric_std.all;
library ocpi; use ocpi.types.all; -- remove this to avoid all ocpi name collisions
architecture rtl of bias_vhdl1_worker is
begin
end rtl;
