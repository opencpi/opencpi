../../../sobel_32f.rcc/target-linux-c6-x86_64/generics.vhd