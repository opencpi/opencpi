../../../bias_param.rcc/target-1-macos-10_9-x86_64/generics.vhd