-- THIS FILE WAS ORIGINALLY GENERATED ON Sun Sep 13 08:43:35 2015 EDT
-- BASED ON THE FILE: cstest.xml
-- YOU *ARE* EXPECTED TO EDIT IT
-- This file initially contains the architecture skeleton for worker: cstest

library IEEE; use IEEE.std_logic_1164.all; use ieee.numeric_std.all;
library ocpi; use ocpi.types.all; -- remove this to avoid all ocpi name collisions
architecture rtl of cstest_worker is
begin
  dummy <= '1';
end rtl;
