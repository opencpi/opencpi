../../../bias_param.rcc/target-2-macos-10_9-x86_64/generics.vhd