../../../convert_s16_f32.rcc/target-linux-c6-x86_64/generics.vhd