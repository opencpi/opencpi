-- THIS FILE WAS ORIGINALLY GENERATED ON Fri Sep 28 22:32:32 2012 EDT
-- BASED ON THE FILE: gen/sym_fir_real.xml
-- YOU *ARE* EXPECTED TO EDIT IT
-- This file initially contains the architecture skeleton for worker: sym_fir_real

library IEEE; use IEEE.std_logic_1164.all; use ieee.numeric_std.all;
library ocpi; use ocpi.types.all; -- remove this to avoid all ocpi name collisions
architecture rtl of sym_fir_real_worker is
begin
end rtl;
