../../../sym_fir_real.rcc/target-linux-c6-x86_64/generics.vhd