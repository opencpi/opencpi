../../../splitter2x2.rcc/target-linux-c6-x86_64/generics.vhd