// THIS FILE WAS ORIGINALLY GENERATED ON Thu Sep 20 16:25:26 2012 EDT
// BASED ON THE FILE: mixer_complex.xml
// YOU ARE EXPECTED TO EDIT IT
// This file contains the implementation skeleton for worker: mixer_complex

`include "mixer_complex-impl.vh"



endmodule //mixer_complex
