// THIS FILE WAS ORIGINALLY GENERATED ON Thu Sep 20 16:14:53 2012 EDT
// BASED ON THE FILE: dsample_complex.xml
// YOU ARE EXPECTED TO EDIT IT
// This file contains the implementation skeleton for worker: dsample_complex

`include "dsample_complex-impl.vh"



endmodule //dsample_complex
