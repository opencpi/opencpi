-- THIS FILE WAS ORIGINALLY GENERATED ON Mon Jun  3 17:13:21 2013 EDT
-- BASED ON THE FILE: gen/file_write.xml
-- YOU *ARE* EXPECTED TO EDIT IT
-- This file initially contains the architecture skeleton for worker: file_write

library IEEE; use IEEE.std_logic_1164.all; use ieee.numeric_std.all;
library ocpi; use ocpi.types.all; -- remove this to avoid all ocpi name collisions
architecture rtl of file_write_worker is
begin
end rtl;
