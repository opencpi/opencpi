// THIS FILE WAS ORIGINALLY GENERATED ON Thu Sep 20 16:24:11 2012 EDT
// BASED ON THE FILE: dds_complex.xml
// YOU ARE EXPECTED TO EDIT IT
// This file contains the implementation skeleton for worker: dds_complex

`include "dds_complex-impl.vh"



endmodule //dds_complex
