/*
 * This file is protected by Copyright. Please refer to the COPYRIGHT file
 * distributed with this source distribution.
 *
 * This file is part of OpenCPI <http://www.opencpi.org>
 *
 * OpenCPI is free software: you can redistribute it and/or modify it under the
 * terms of the GNU Lesser General Public License as published by the Free
 * Software Foundation, either version 3 of the License, or (at your option) any
 * later version.
 *
 * OpenCPI is distributed in the hope that it will be useful, but WITHOUT ANY
 * WARRANTY; without even the implied warranty of MERCHANTABILITY or FITNESS FOR
 * A PARTICULAR PURPOSE. See the GNU Lesser General Public License for more
 * details.
 *
 * You should have received a copy of the GNU Lesser General Public License
 * along with this program. If not, see <http://www.gnu.org/licenses/>.
 */

localparam OCPI_OCP_MCMD_WRITE = 3'h1;
localparam OCPI_OCP_MCMD_READ  = 3'h2;
localparam OCPI_OCP_MCMD_IDLE  = 3'h0;
localparam OCPI_OCP_SRESP_NULL = 2'h0;
localparam OCPI_OCP_SRESP_DVA  = 2'h1;
localparam OCPI_OCP_SRESP_FAIL = 2'h2;
localparam OCPI_OCP_SRESP_ERR  = 2'h3;


