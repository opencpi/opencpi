../../../../assets/hdl/devices/ad9361_config.hdl/signals.vhd