../../../min_eigen_val.rcc/target-linux-c6-x86_64/generics.vhd