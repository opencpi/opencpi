../../../corner_eigen_vals_vecs.rcc/target-macos-10_9-x86_64/generics.vhd