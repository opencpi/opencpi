-- This file is protected by Copyright. Please refer to the COPYRIGHT file
-- distributed with this source distribution.
--
-- This file is part of OpenCPI <http:--www.opencpi.org>
--
-- OpenCPI is free software: you can redistribute it and/or modify it under the
-- terms of the GNU Lesser General Public License as published by the Free
-- Software Foundation, either version 3 of the License, or (at your option) any
-- later version.
--
-- OpenCPI is distributed in the hope that it will be useful, but WITHOUT ANY
-- WARRANTY; without even the implied warranty of MERCHANTABILITY or FITNESS FOR
-- A PARTICULAR PURPOSE. See the GNU Lesser General Public License for more
-- details.
--
-- You should have received a copy of the GNU Lesser General Public License
-- along with this program. If not, see <http:--www.gnu.org/licenses/>.

-- This file is our wrapper around the processing_system8 IP as generated by
-- ps8.tcl.
-- There is no logic here, just providing a simpler interface for the platform worker
-- that uses it.
library IEEE; use IEEE.std_logic_1164.all; use ieee.numeric_std.all;
library ocpi; use ocpi.types.all; -- remove this to avoid all ocpi name collisions
library zynq_ultra; use zynq_ultra.zynq_ultra_pkg.all;
library axi; use axi.axi_pkg.all;
entity zynq_ultra_ps_e is
  port(
    ps_in        : in    pl2ps_t;
    ps_out       : out   ps2pl_t;
    m_axi_hp_in  : in    m_axi_hp_in_array_t(0 to C_M_AXI_HP_COUNT-1);
    m_axi_hp_out : out   m_axi_hp_out_array_t(0 to C_M_AXI_HP_COUNT-1);
    s_axi_hp_in  : in    s_axi_hp_in_array_t(0 to C_S_AXI_HP_COUNT-1);
    s_axi_hp_out : out   s_axi_hp_out_array_t(0 to C_S_AXI_HP_COUNT-1)
    );
end entity zynq_ultra_ps_e;
architecture rtl of zynq_ultra_ps_e is
  -- Various SLV arrays of different SLV widths for use below
  type vec_49_array_t is array (natural range <>) of std_logic_vector(48 downto 0);
  type vec_40_array_t is array (natural range <>) of std_logic_vector(39 downto 0);
  type vec_32_array_t is array (natural range <>) of std_logic_vector(31 downto 0);
  type vec_16_array_t is array (natural range <>) of std_logic_vector(15 downto 0);
  type vec_8_array_t is array (natural range <>) of std_logic_vector(7 downto 0);
  type vec_6_array_t is array (natural range <>) of std_logic_vector(5 downto 0);
  type vec_4_array_t is array (natural range <>) of std_logic_vector(3 downto 0);

  -- Some AXI signals have bit-width mismatches between the UltraScale PS8 and
  -- the OpenCPI AXI primitive. These intermediate signals below are used to
  -- compensate for the mismatches by leaving higher-order unused signals open
  -- or tied to '0'
  signal maxigp_awids   : vec_16_array_t(0 to C_M_AXI_HP_COUNT-1);
  signal maxigp_awaddrs : vec_40_array_t(0 to C_M_AXI_HP_COUNT-1);
  signal maxigp_awlens  : vec_8_array_t (0 to C_M_AXI_HP_COUNT-1);

  signal maxigp_arids   : vec_16_array_t(0 to C_M_AXI_HP_COUNT-1);
  signal maxigp_araddrs : vec_40_array_t(0 to C_M_AXI_HP_COUNT-1);
  signal maxigp_arlens  : vec_8_array_t (0 to C_M_AXI_HP_COUNT-1);

  signal maxigp_bids    : vec_16_array_t(0 to C_M_AXI_HP_COUNT-1);
  signal maxigp_rids    : vec_16_array_t(0 to C_M_AXI_HP_COUNT-1);

  signal saxigp_awaddrs : vec_49_array_t(0 to C_S_AXI_HP_COUNT-1);
  signal saxigp_awlens  : vec_8_array_t (0 to C_S_AXI_HP_COUNT-1);

  signal saxigp_araddrs : vec_49_array_t(0 to C_S_AXI_HP_COUNT-1);
  signal saxigp_arlens  : vec_8_array_t (0 to C_S_AXI_HP_COUNT-1);

  signal saxigp_racounts : vec_4_array_t(0 to C_S_AXI_HP_COUNT-1);
  signal saxigp_wacounts : vec_4_array_t(0 to C_S_AXI_HP_COUNT-1);

begin

  -- tie higher-order unused signals to '0' and connect only needed ones
  m : for i in 0 to C_M_AXI_HP_COUNT-1 generate
    m_axi_hp_out(i).AW.ID <= maxigp_awids(i)(11 downto 0);
    m_axi_hp_out(i).AR.ID <= maxigp_arids(i)(11 downto 0);
    m_axi_hp_out(i).AW.LOCK(1) <= '0';
    m_axi_hp_out(i).AW.ISSUECAP1_EN <= '0';
    m_axi_hp_out(i).AR.ISSUECAP1_EN <= '0';
    maxigp_bids(i)(11 downto 0)  <= m_axi_hp_in(0).B.ID;
    maxigp_bids(i)(15 downto 12) <= (others =>'0');
    maxigp_rids(i)(11 downto 0) <= m_axi_hp_in(0).R.ID;
    maxigp_rids(i)(15 downto 12) <= (others =>'0');
  end generate;

  s : for i in 0 to C_S_AXI_HP_COUNT-1 generate
    s_axi_hp_out(i).AR.COUNT <= saxigp_racounts(i)(2 downto 0);
    s_axi_hp_out(i).AW.COUNT(5 downto 4) <= (others => '0');
    saxigp_awaddrs(i)(31 downto 0)  <= s_axi_hp_in(0).AW.ADDR;
    saxigp_awaddrs(i)(48 downto 32) <= (others =>'0');
    saxigp_araddrs(i)(31 downto 0)  <= s_axi_hp_in(0).AR.ADDR;
    saxigp_araddrs(i)(48 downto 32) <= (others =>'0');
    saxigp_awlens(i)(3 downto 0)  <= s_axi_hp_in(0).AW.LEN;
    saxigp_awlens(i)(7 downto 4) <= (others =>'0');
    saxigp_arlens(i)(3 downto 0)  <= s_axi_hp_in(0).AR.LEN;
    saxigp_arlens(i)(7 downto 4) <= (others =>'0');
  end generate;

  -- Connect the Verilog PS8 wrapper to the VHDL axi records to abstract the interface
  ps : zynq_ultra_ps_e_v3_2_1_zynq_ultra_ps_e
    generic map(
      C_MAXIGP0_DATA_WIDTH => 32,
      C_MAXIGP1_DATA_WIDTH => 32,
      C_MAXIGP2_DATA_WIDTH => 128,

      C_SAXIGP0_DATA_WIDTH => 128,
      C_SAXIGP1_DATA_WIDTH => 128,
      C_SAXIGP2_DATA_WIDTH => 64,
      C_SAXIGP3_DATA_WIDTH => 64,
      C_SAXIGP4_DATA_WIDTH => 64,
      C_SAXIGP5_DATA_WIDTH => 64,
      C_SAXIGP6_DATA_WIDTH => 128,
      C_SD0_INTERNAL_BUS_WIDTH => 8,
      C_SD1_INTERNAL_BUS_WIDTH => 8,
      C_PL_CLK0_BUF => "FALSE", -- was TRUE in default
      C_PL_CLK1_BUF => "FALSE", -- was TRUE in default -- FALSE in TRD
      C_PL_CLK2_BUF => "FALSE", -- was TRUE in default -- FALSE in TRD
      C_PL_CLK3_BUF => "FALSE", -- was TRUE in default -- FALSE in TRD

      C_NUM_F2P_0_INTR_INPUTS => 0,  -- 1 in TRD
      C_NUM_F2P_1_INTR_INPUTS => 0,  -- 1 in TRD

      C_NUM_FABRIC_RESETS => 1,
      C_EMIO_GPIO_WIDTH => 60, -- 95 in TRD

      -- C_TRISTATE_INVERTED => 1,

      C_USE_DIFF_RW_CLK_GP0 => 0,
      C_USE_DIFF_RW_CLK_GP1 => 0,
      C_USE_DIFF_RW_CLK_GP2 => 0,
      C_USE_DIFF_RW_CLK_GP3 => 0,
      C_USE_DIFF_RW_CLK_GP4 => 0,
      C_USE_DIFF_RW_CLK_GP5 => 0,
      C_USE_DIFF_RW_CLK_GP6 => 0,

      C_TRACE_PIPELINE_WIDTH => 8,
      C_EN_EMIO_TRACE => 0,
      C_EN_FIFO_ENET0 => 0,
      C_EN_FIFO_ENET1 => 0,
      C_EN_FIFO_ENET2 => 0,
      C_EN_FIFO_ENET3 => 0,
      C_TRACE_DATA_WIDTH => 32,

      C_USE_DEBUG_TEST => 0,
      C_DP_USE_AUDIO => 0,
      C_DP_USE_VIDEO => 0 -- 1 in TRD
    )
    port map(
-- maxigp0
      maxihpm0_fpd_aclk => m_axi_hp_in(0).ACLK,
      dp_video_ref_clk => open,
      dp_audio_ref_clk => open,
      maxigp0_awid => maxigp_awids(0), --[15:0]
      maxigp0_awaddr => maxigp_awaddrs(0), --[39:0]
      maxigp0_awlen => maxigp_awlens(0), --[7:0]
      maxigp0_awsize => m_axi_hp_out(0).AW.SIZE, --[2:0]
      maxigp0_awburst => m_axi_hp_out(0).AW.BURST, --[1:0]
      maxigp0_awlock => m_axi_hp_out(0).AW.LOCK(0),
      maxigp0_awcache => m_axi_hp_out(0).AW.CACHE, --[3:0]
      maxigp0_awprot => m_axi_hp_out(0).AW.PROT, --[2:0]
      maxigp0_awvalid => m_axi_hp_out(0).AW.VALID,
      maxigp0_awuser => open, --[15:0]
      maxigp0_awready => m_axi_hp_in(0).AW.READY,
      maxigp0_wdata => m_axi_hp_out(0).W.DATA, --[C_MAXIGP0_DATA_WIDTH-1 :0]
      maxigp0_wstrb => m_axi_hp_out(0).W.STRB, --[(C_MAXIGP0_DATA_WIDTH/8)-1 :0]
      maxigp0_wlast => m_axi_hp_out(0).W.LAST,
      maxigp0_wvalid => m_axi_hp_out(0).W.VALID,
      maxigp0_wready => m_axi_hp_in(0).W.READY,
      maxigp0_bid => maxigp_bids(0), --[15:0]
      maxigp0_bresp => m_axi_hp_in(0).B.RESP, --[1:0]
      maxigp0_bvalid => m_axi_hp_in(0).B.VALID,
      maxigp0_bready => m_axi_hp_out(0).B.READY,
      maxigp0_arid => maxigp_arids(0), --[15:0]
      maxigp0_araddr => maxigp_araddrs(0), --[39:0]
      maxigp0_arlen => maxigp_arlens(0), --[7:0]
      maxigp0_arsize => m_axi_hp_out(0).AR.SIZE, --[2:0]
      maxigp0_arburst => m_axi_hp_out(0).AR.BURST, --[1:0]
      maxigp0_arlock => m_axi_hp_out(0).AR.LOCK(0),
      maxigp0_arcache => m_axi_hp_out(0).AR.CACHE, --[3:0]
      maxigp0_arprot => m_axi_hp_out(0).AR.PROT, --[2:0]
      maxigp0_arvalid => m_axi_hp_out(0).AR.VALID,
      maxigp0_aruser => open, --[15:0]
      maxigp0_arready => m_axi_hp_in(0).AR.READY,
      maxigp0_rid => maxigp_rids(0), --[15:0]
      maxigp0_rdata => m_axi_hp_in(0).R.DATA, --[C_MAXIGP0_DATA_WIDTH-1 :0]
      maxigp0_rresp => m_axi_hp_in(0).R.RESP, --[1:0]
      maxigp0_rlast => m_axi_hp_in(0).R.LAST,
      maxigp0_rvalid => m_axi_hp_in(0).R.VALID,
      maxigp0_rready => m_axi_hp_out(0).R.READY,
      maxigp0_awqos => m_axi_hp_out(0).AW.QOS, --[3:0]
      maxigp0_arqos => m_axi_hp_out(0).AR.QOS, --[3:0]

-- maxigp1
      maxihpm1_fpd_aclk => m_axi_hp_in(1).ACLK,
      maxigp1_awid => maxigp_awids(1),
      maxigp1_awaddr => maxigp_awaddrs(1),
      maxigp1_awlen => maxigp_awlens(1),
      maxigp1_awsize => m_axi_hp_out(1).AW.SIZE, --[2:0]
      maxigp1_awburst => m_axi_hp_out(1).AW.BURST, --[1:0]
      maxigp1_awlock => m_axi_hp_out(1).AW.LOCK(0),
      maxigp1_awcache => m_axi_hp_out(1).AW.CACHE, --[3:0]
      maxigp1_awprot => m_axi_hp_out(1).AW.PROT, --[2:0]
      maxigp1_awvalid => m_axi_hp_out(1).AW.VALID,
      maxigp1_awuser => open, --[15:0]
      maxigp1_awready => m_axi_hp_in(1).AW.READY,
      maxigp1_wdata => m_axi_hp_out(1).W.DATA, --[C_MAXIGP1_DATA_WIDTH-1 :0]
      maxigp1_wstrb => m_axi_hp_out(1).W.STRB, --[(C_MAXIGP1_DATA_WIDTH/8)-1 :0]
      maxigp1_wlast => m_axi_hp_out(1).W.LAST,
      maxigp1_wvalid => m_axi_hp_out(1).W.VALID,
      maxigp1_wready => m_axi_hp_in(1).W.READY,
      maxigp1_bid => maxigp_bids(1), --m_axi_hp_in(1).B.ID, --[15:0]
      maxigp1_bresp => m_axi_hp_in(1).B.RESP, --[1:0]
      maxigp1_bvalid => m_axi_hp_in(1).B.VALID,
      maxigp1_bready => m_axi_hp_out(1).B.READY,
      maxigp1_arid => maxigp_arids(1),
      maxigp1_araddr => maxigp_araddrs(1),
      maxigp1_arlen => maxigp_arlens(1),
      maxigp1_arsize => m_axi_hp_out(1).AR.SIZE, --[2:0]
      maxigp1_arburst => m_axi_hp_out(1).AR.BURST, --[1:0]
      maxigp1_arlock => m_axi_hp_out(1).AR.LOCK(0),
      maxigp1_arprot => m_axi_hp_out(1).AR.PROT, --[2:0]
      maxigp1_arcache => m_axi_hp_out(1).AR.CACHE, --[3:0]
      maxigp1_arvalid => m_axi_hp_out(1).AR.VALID,
      maxigp1_aruser => open, --[15:0]
      maxigp1_arready => m_axi_hp_in(1).AR.READY,
      maxigp1_rid => maxigp_rids(1), --[15:0]
      maxigp1_rdata => m_axi_hp_in(1).R.DATA, --[C_MAXIGP1_DATA_WIDTH-1 :0]
      maxigp1_rresp => m_axi_hp_in(1).R.RESP, --[1:0]
      maxigp1_rlast => m_axi_hp_in(1).R.LAST,
      maxigp1_rvalid => m_axi_hp_in(1).R.VALID,
      maxigp1_rready => m_axi_hp_out(1).R.READY,
      maxigp1_awqos => m_axi_hp_out(1).AW.QOS, --[3:0]
      maxigp1_arqos => m_axi_hp_out(1).AR.QOS, --[3:0]
-- maxigp2
      -- NOT USING
      maxihpm0_lpd_aclk => '0',
      maxigp2_awid => open, -- m_axi_hp_out(2).AW.ID, --[15:0]
      maxigp2_awaddr => open, -- m_axi_hp_out(2).AW.ADDR, --[39:0]
      maxigp2_awlen => open, -- m_axi_hp_out(2).AW.LEN, --[7:0]
      maxigp2_awsize => open, -- m_axi_hp_out(2).AW.SIZE, --[2:0]
      maxigp2_awburst => open, -- m_axi_hp_out(2).AW.BURST, --[1:0]
      maxigp2_awlock => open, -- m_axi_hp_out(2).AW.LOCK(0),
      maxigp2_awcache => open, -- m_axi_hp_out(2).AW.CACHE, --[3:0]
      maxigp2_awprot => open, -- m_axi_hp_out(2).AW.PROT, --[2:0]
      maxigp2_awvalid => open, -- m_axi_hp_out(2).AW.VALID,
      maxigp2_awuser => open, -- m_axi_hp_out(2).AWUSER, --[15:0]
      maxigp2_awready => '0', -- m_axi_hp_in(2).AW.READY,
      maxigp2_wdata => open, -- m_axi_hp_out(2).W.DATA, --[C_MAXIGP2_DATA_WIDTH-1 :0]
      maxigp2_wstrb => open, -- m_axi_hp_out(2).W.STRB, --[(C_MAXIGP2_DATA_WIDTH/8)-1 :0]
      maxigp2_wlast => open, -- m_axi_hp_out(2).W.LAST,
      maxigp2_wvalid => open, -- m_axi_hp_out(2).W.VALID,
      maxigp2_wready => '0', -- m_axi_hp_in(2).W.READY,
      maxigp2_bid => (others => '0'), -- m_axi_hp_in(2).B.ID, --[15:0]
      maxigp2_bresp => (others => '0'), -- m_axi_hp_in(2).B.RESP, --[1:0]
      maxigp2_bvalid => '0', -- m_axi_hp_in(2).B.VALID,
      maxigp2_bready => open, -- m_axi_hp_out(2).B.READY,
      maxigp2_arid => open, -- m_axi_hp_out(2).AR.ID, --[15:0]
      maxigp2_araddr => open, -- m_axi_hp_out(2).AR.ADDR, --[39:0]
      maxigp2_arlen => open, -- m_axi_hp_out(2).AR.LEN, --[7:0]
      maxigp2_arsize => open, -- m_axi_hp_out(2).AR.SIZE, --[2:0]
      maxigp2_arburst => open, -- m_axi_hp_out(2).AR.BURST, --[1:0]
      maxigp2_arlock => open, -- m_axi_hp_out(2).AR.LOCK(0),
      maxigp2_arcache => open, -- m_axi_hp_out(2).AR.CACHE, --[3:0]
      maxigp2_arprot => open, -- m_axi_hp_out(2).AR.PROT, --[2:0]
      maxigp2_arvalid => open, -- m_axi_hp_out(2).AR.VALID,
      maxigp2_aruser => open, -- m_axi_hp_out(2).ARUSER, --[15:0]
      maxigp2_arready => '0', -- m_axi_hp_in(2).AR.READY,
      maxigp2_rid => (others => '0'), -- m_axi_hp_in(2).R.ID, --[15:0]
      maxigp2_rdata => (others => '0'), -- m_axi_hp_in(2).R.DATA, --[C_MAXIGP2_DATA_WIDTH-1 :0]
      maxigp2_rresp => (others => '0'), -- m_axi_hp_in(2).R.RESP, --[1:0]
      maxigp2_rlast => '0', -- m_axi_hp_in(2).R.LAST,
      maxigp2_rvalid => '0', -- m_axi_hp_in(2).R.VALID,
      maxigp2_rready => open, -- m_axi_hp_out(2).R.READY,
      maxigp2_awqos => open, -- m_axi_hp_out(2).AW.QOS, --[3:0]
      maxigp2_arqos => open, -- m_axi_hp_out(2).AR.QOS, --[3:0]
-- saxigp0
      -- NOT USING
      saxihpc0_fpd_aclk => '0', -- saxihpc0_fpd_aclk => s_axi_hp_in(0).ACLK,
      saxihpc0_fpd_rclk => '0',
      saxihpc0_fpd_wclk => '0',
      saxigp0_aruser => '0', -- s_axi_hp_in(0).ARUSER,
      saxigp0_awuser => '0', -- s_axi_hp_in(0).AWUSER,
      saxigp0_awid => (others => '0'), -- s_axi_hp_in(0).AW.ID, --[5:0]
      saxigp0_awaddr => (others => '0'), -- s_axi_hp_in(0).AW.ADDR, --[48:0]
      saxigp0_awlen => (others => '0'), -- s_axi_hp_in(0).AW.LEN, --[7:0]
      saxigp0_awsize => (others => '0'), -- s_axi_hp_in(0).AW.SIZE, --[2:0]
      saxigp0_awburst => (others => '0'), -- s_axi_hp_in(0).AW.BURST, --[1:0]
      saxigp0_awlock => '0', -- s_axi_hp_in(0).AW.LOCK(0),
      saxigp0_awcache => (others => '0'), -- s_axi_hp_in(0).AW.CACHE, --[3:0]
      saxigp0_awprot => (others => '0'), -- s_axi_hp_in(0).AW.PROT, --[2:0]
      saxigp0_awvalid => '0', -- s_axi_hp_in(0).AW.VALID,
      saxigp0_awready => open, -- s_axi_hp_out(0).AW.READY,
      saxigp0_wdata => (others => '0'), -- s_axi_hp_in(0).W.DATA, --[C_SAXIGP0_DATA_WIDTH-1:0]
      saxigp0_wstrb => (others => '0'), -- s_axi_hp_in(0).W.STRB, --[(C_SAXIGP0_DATA_WIDTH/8) -1 :0]
      saxigp0_wlast => '0', -- s_axi_hp_in(0).W.LAST,
      saxigp0_wvalid => '0', -- s_axi_hp_in(0).W.VALID,
      saxigp0_wready => open, -- s_axi_hp_out(0).W.READY,
      saxigp0_bid => open, -- s_axi_hp_out(0).B.ID, --[5:0]
      saxigp0_bresp => open, -- s_axi_hp_out(0).B.RESP, --[1:0]
      saxigp0_bvalid => open, -- s_axi_hp_out(0).B.VALID,
      saxigp0_bready => '0', -- s_axi_hp_in(0).B.READY,
      saxigp0_arid => (others => '0'), -- s_axi_hp_in(0).AR.ID, --[5:0]
      saxigp0_araddr => (others => '0'), -- s_axi_hp_in(0).AR.ADDR, --[48:0]
      saxigp0_arlen => (others => '0'), -- s_axi_hp_in(0).AR.LEN, --[7:0]
      saxigp0_arsize => (others => '0'), -- s_axi_hp_in(0).AR.SIZE, --[2:0]
      saxigp0_arburst => (others => '0'), -- s_axi_hp_in(0).AR.BURST, --[1:0]
      saxigp0_arlock => '0', -- s_axi_hp_in(0).AR.LOCK(0),
      saxigp0_arcache => (others => '0'), -- s_axi_hp_in(0).AR.CACHE, --[3:0]
      saxigp0_arprot => (others => '0'), -- s_axi_hp_in(0).AR.PROT, --[2:0]
      saxigp0_arvalid => '0', -- s_axi_hp_in(0).AR.VALID,
      saxigp0_arready => open, -- s_axi_hp_out(0).AR.READY,
      saxigp0_rid => open, -- s_axi_hp_out(0).R.ID, --[5:0]
      saxigp0_rdata => open, -- s_axi_hp_out(0).R.DATA, --[C_SAXIGP0_DATA_WIDTH-1:0]
      saxigp0_rresp => open, -- s_axi_hp_out(0).R.RESP, --[1:0]
      saxigp0_rlast => open, -- s_axi_hp_out(0).R.LAST,
      saxigp0_rvalid => open, -- s_axi_hp_out(0).R.VALID,
      saxigp0_rready => '0', -- s_axi_hp_in(0).R.READY,
      saxigp0_awqos => (others => '0'), -- s_axi_hp_in(0).AW.QOS, --[3:0]
      saxigp0_arqos => (others => '0'), -- s_axi_hp_in(0).AR.QOS, --[3:0]
      saxigp0_rcount => open, -- s_axi_hp_out(0).R.COUNT, --[7:0]
      saxigp0_wcount => open, -- s_axi_hp_out(0).W.COUNT, --[7:0]
      saxigp0_racount => open, -- s_axi_hp_out(0).AR.COUNT, --[3:0]
      saxigp0_wacount => open, -- s_axi_hp_out(0).AW.COUNT, --[3:0]
-- saxigp1
      -- NOT USING
      saxihpc1_fpd_aclk => '0', -- s_axi_hp_in(1).ACLK,
      saxihpc1_fpd_rclk => '0',
      saxihpc1_fpd_wclk => '0',
      saxigp1_aruser => '0', -- s_axi_hp_in(1).ARUSER,
      saxigp1_awuser => '0', -- s_axi_hp_in(1).AWUSER,
      saxigp1_awid => (others => '0'), -- s_axi_hp_in(1).AW.ID, --[5:0]
      saxigp1_awaddr => (others => '0'), -- s_axi_hp_in(1).AW.ADDR, --[48:0]
      saxigp1_awlen => (others => '0'), -- s_axi_hp_in(1).AW.LEN, --[7:0]
      saxigp1_awsize => (others => '0'), -- s_axi_hp_in(1).AW.SIZE, --[2:0]
      saxigp1_awburst => (others => '0'), -- s_axi_hp_in(1).AW.BURST, --[1:0]
      saxigp1_awlock => '0', -- s_axi_hp_in(1).AW.LOCK(0),
      saxigp1_awcache => (others => '0'), -- s_axi_hp_in(1).AW.CACHE, --[3:0]
      saxigp1_awprot => (others => '0'), -- s_axi_hp_in(1).AW.PROT, --[2:0]
      saxigp1_awvalid => '0', -- s_axi_hp_in(1).AW.VALID,
      saxigp1_awready => open, -- s_axi_hp_out(1).AW.READY,
      saxigp1_wdata => (others => '0'), -- s_axi_hp_in(1).W.DATA, --[C_SAXIGP1_DATA_WIDTH-1:0]
      saxigp1_wstrb => (others => '0'), -- s_axi_hp_in(1).W.STRB, --[(C_SAXIGP1_DATA_WIDTH/8) -1 :0]
      saxigp1_wlast => '0', -- s_axi_hp_in(1).W.LAST,
      saxigp1_wvalid => '0', -- s_axi_hp_in(1).W.VALID,
      saxigp1_wready => open, -- s_axi_hp_out(1).W.READY,
      saxigp1_bid => open, -- s_axi_hp_out(1).B.ID, --[5:0]
      saxigp1_bresp => open, -- s_axi_hp_out(1).B.RESP, --[1:0]
      saxigp1_bvalid => open, -- s_axi_hp_out(1).B.VALID,
      saxigp1_bready => '0', -- s_axi_hp_in(1).B.READY,
      saxigp1_arid => (others => '0'), -- s_axi_hp_in(1).AR.ID, --[5:0]
      saxigp1_araddr => (others => '0'), -- s_axi_hp_in(1).AR.ADDR, --[48:0]
      saxigp1_arlen => (others => '0'), -- s_axi_hp_in(1).AR.LEN, --[7:0]
      saxigp1_arsize => (others => '0'), -- s_axi_hp_in(1).AR.SIZE, --[2:0]
      saxigp1_arburst => (others => '0'), -- s_axi_hp_in(1).AR.BURST, --[1:0]
      saxigp1_arlock => '0', -- s_axi_hp_in(1).AR.LOCK(0),
      saxigp1_arcache => (others => '0'), -- s_axi_hp_in(1).AR.CACHE, --[3:0]
      saxigp1_arprot => (others => '0'), -- s_axi_hp_in(1).AR.PROT, --[2:0]
      saxigp1_arvalid => '0', -- s_axi_hp_in(1).AR.VALID,
      saxigp1_arready => open, -- s_axi_hp_out(1).AR.READY,
      saxigp1_rid => open, -- s_axi_hp_out(1).R.ID, --[5:0]
      saxigp1_rdata => open, -- s_axi_hp_out(1).R.DATA, --[C_SAXIGP1_DATA_WIDTH-1:0]
      saxigp1_rresp => open, -- s_axi_hp_out(1).R.RESP, --[1:0]
      saxigp1_rlast => open, -- s_axi_hp_out(1).R.LAST,
      saxigp1_rvalid => open, -- s_axi_hp_out(1).R.VALID,
      saxigp1_rready => '0', -- s_axi_hp_in(1).R.READY,
      saxigp1_awqos => (others => '0'), -- s_axi_hp_in(1).AW.QOS, --[3:0]
      saxigp1_arqos => (others => '0'), -- s_axi_hp_in(1).AR.QOS, --[3:0]
      saxigp1_rcount => open, -- s_axi_hp_out(1).R.COUNT, --[7:0]
      saxigp1_wcount => open, -- s_axi_hp_out(1).W.COUNT, --[7:0]
      saxigp1_racount => open, -- s_axi_hp_out(1).AR.COUNT, --[3:0]
      saxigp1_wacount => open, -- s_axi_hp_out(1).AW.COUNT, --[3:0]
-- saxigp2
      saxihp0_fpd_aclk => s_axi_hp_in(0).ACLK,
      saxihp0_fpd_rclk => '0',
      saxihp0_fpd_wclk => '0',
      saxigp2_aruser => '0',
      saxigp2_awuser => '0',
      saxigp2_awid => s_axi_hp_in(0).AW.ID(5 downto 0), --[5:0]
      saxigp2_awaddr => saxigp_awaddrs(0), --[48:0]
      saxigp2_awlen => saxigp_awlens(0), --[7:0]
      saxigp2_awsize => s_axi_hp_in(0).AW.SIZE, --[2:0]
      saxigp2_awburst => s_axi_hp_in(0).AW.BURST, --[1:0]
      saxigp2_awlock => s_axi_hp_in(0).AW.LOCK(0),
      saxigp2_awcache => s_axi_hp_in(0).AW.CACHE, --[3:0]
      saxigp2_awprot => s_axi_hp_in(0).AW.PROT, --[2:0]
      saxigp2_awvalid => s_axi_hp_in(0).AW.VALID,
      saxigp2_awready => s_axi_hp_out(0).AW.READY,
      saxigp2_wdata => s_axi_hp_in(0).W.DATA, --[C_SAXIGP2_DATA_WIDTH-1:0]
      saxigp2_wstrb => s_axi_hp_in(0).W.STRB, --[(C_SAXIGP2_DATA_WIDTH/8) -1 :0]
      saxigp2_wlast => s_axi_hp_in(0).W.LAST,
      saxigp2_wvalid => s_axi_hp_in(0).W.VALID,
      saxigp2_wready => s_axi_hp_out(0).W.READY,
      saxigp2_bid => s_axi_hp_out(0).B.ID(5 downto 0), --[5:0]
      saxigp2_bresp => s_axi_hp_out(0).B.RESP, --[1:0]
      saxigp2_bvalid => s_axi_hp_out(0).B.VALID,
      saxigp2_bready => s_axi_hp_in(0).B.READY,
      saxigp2_arid => s_axi_hp_in(0).AR.ID(5 downto 0), --[5:0]
      saxigp2_araddr => saxigp_araddrs(0), --[48:0]
      saxigp2_arlen => saxigp_arlens(0), --[7:0]
      saxigp2_arsize => s_axi_hp_in(0).AR.SIZE, --[2:0]
      saxigp2_arburst => s_axi_hp_in(0).AR.BURST, --[1:0]
      saxigp2_arlock => s_axi_hp_in(0).AR.LOCK(0),
      saxigp2_arcache => s_axi_hp_in(0).AR.CACHE, --[3:0]
      saxigp2_arprot => s_axi_hp_in(0).AR.PROT, --[2:0]
      saxigp2_arvalid => s_axi_hp_in(0).AR.VALID,
      saxigp2_arready => s_axi_hp_out(0).AR.READY,
      saxigp2_rid => s_axi_hp_out(0).R.ID(5 downto 0), --[5:0]
      saxigp2_rdata => s_axi_hp_out(0).R.DATA, --[C_SAXIGP2_DATA_WIDTH-1:0]
      saxigp2_rresp => s_axi_hp_out(0).R.RESP, --[1:0]
      saxigp2_rlast => s_axi_hp_out(0).R.LAST,
      saxigp2_rvalid => s_axi_hp_out(0).R.VALID,
      saxigp2_rready => s_axi_hp_in(0).R.READY,
      saxigp2_awqos => s_axi_hp_in(0).AW.QOS, --[3:0]
      saxigp2_arqos => s_axi_hp_in(0).AR.QOS, --[3:0]
      saxigp2_rcount => s_axi_hp_out(0).R.COUNT, --[7:0]
      saxigp2_wcount => s_axi_hp_out(0).W.COUNT, --[7:0]
      saxigp2_racount => saxigp_racounts(0), --[3:0]
      saxigp2_wacount => s_axi_hp_out(0).AW.COUNT(3 downto 0), --[3:0]
-- saxigp3
      saxihp1_fpd_aclk => s_axi_hp_in(1).ACLK,
      saxihp1_fpd_rclk => '0',
      saxihp1_fpd_wclk => '0',
      saxigp3_aruser => '0',
      saxigp3_awuser => '0',
      saxigp3_awid => s_axi_hp_in(1).AW.ID(5 downto 0), --[5:0]
      saxigp3_awaddr => saxigp_awaddrs(1), --[48:0]
      saxigp3_awlen => saxigp_awlens(1), --[7:0]
      saxigp3_awsize => s_axi_hp_in(1).AW.SIZE, --[2:0]
      saxigp3_awburst => s_axi_hp_in(1).AW.BURST, --[1:0]
      saxigp3_awlock => s_axi_hp_in(1).AW.LOCK(0),
      saxigp3_awcache => s_axi_hp_in(1).AW.CACHE, --[3:0]
      saxigp3_awprot => s_axi_hp_in(1).AW.PROT, --[2:0]
      saxigp3_awvalid => s_axi_hp_in(1).AW.VALID,
      saxigp3_awready => s_axi_hp_out(1).AW.READY,
      saxigp3_wdata => s_axi_hp_in(1).W.DATA, --[C_SAXIGP3_DATA_WIDTH-1:0]
      saxigp3_wstrb => s_axi_hp_in(1).W.STRB, --[(C_SAXIGP3_DATA_WIDTH/8) -1 :0]
      saxigp3_wlast => s_axi_hp_in(1).W.LAST,
      saxigp3_wvalid => s_axi_hp_in(1).W.VALID,
      saxigp3_wready => s_axi_hp_out(1).W.READY,
      saxigp3_bid => s_axi_hp_out(1).B.ID(5 downto 0), --[5:0]
      saxigp3_bresp => s_axi_hp_out(1).B.RESP, --[1:0]
      saxigp3_bvalid => s_axi_hp_out(1).B.VALID,
      saxigp3_bready => s_axi_hp_in(1).B.READY,
      saxigp3_arid => s_axi_hp_in(1).AR.ID(5 downto 0), --[5:0]
      saxigp3_araddr => saxigp_araddrs(1), --[48:0]
      saxigp3_arlen => saxigp_arlens(1), --[7:0]
      saxigp3_arsize => s_axi_hp_in(1).AR.SIZE, --[2:0]
      saxigp3_arburst => s_axi_hp_in(1).AR.BURST, --[1:0]
      saxigp3_arlock => s_axi_hp_in(1).AR.LOCK(0),
      saxigp3_arcache => s_axi_hp_in(1).AR.CACHE, --[3:0]
      saxigp3_arprot => s_axi_hp_in(1).AR.PROT, --[2:0]
      saxigp3_arvalid => s_axi_hp_in(1).AR.VALID,
      saxigp3_arready => s_axi_hp_out(1).AR.READY,
      saxigp3_rid => s_axi_hp_out(1).R.ID(5 downto 0), --[5:0]
      saxigp3_rdata => s_axi_hp_out(1).R.DATA, --[C_SAXIGP3_DATA_WIDTH-1:0]
      saxigp3_rresp => s_axi_hp_out(1).R.RESP, --[1:0]
      saxigp3_rlast => s_axi_hp_out(1).R.LAST,
      saxigp3_rvalid => s_axi_hp_out(1).R.VALID,
      saxigp3_rready => s_axi_hp_in(1).R.READY,
      saxigp3_awqos => s_axi_hp_in(1).AW.QOS, --[3:0]
      saxigp3_arqos => s_axi_hp_in(1).AR.QOS, --[3:0]
      saxigp3_rcount => s_axi_hp_out(1).R.COUNT, --[7:0]
      saxigp3_wcount => s_axi_hp_out(1).W.COUNT, --[7:0]
      saxigp3_racount => saxigp_racounts(1), --[3:0]
      saxigp3_wacount => s_axi_hp_out(1).AW.COUNT(3 downto 0), --[3:0]
-- saxigp4
      saxihp2_fpd_aclk => s_axi_hp_in(2).ACLK,
      saxihp2_fpd_rclk => '0',
      saxihp2_fpd_wclk => '0',
      saxigp4_aruser => '0',
      saxigp4_awuser => '0',
      saxigp4_awid => s_axi_hp_in(2).AW.ID(5 downto 0), --[5:0]
      saxigp4_awaddr => saxigp_awaddrs(2), --[48:0]
      saxigp4_awlen => saxigp_awlens(2), --[7:0]
      saxigp4_awsize => s_axi_hp_in(2).AW.SIZE, --[2:0]
      saxigp4_awburst => s_axi_hp_in(2).AW.BURST, --[1:0]
      saxigp4_awlock => s_axi_hp_in(2).AW.LOCK(0),
      saxigp4_awcache => s_axi_hp_in(2).AW.CACHE, --[3:0]
      saxigp4_awprot => s_axi_hp_in(2).AW.PROT, --[2:0]
      saxigp4_awvalid => s_axi_hp_in(2).AW.VALID,
      saxigp4_awready => s_axi_hp_out(2).AW.READY,
      saxigp4_wdata => s_axi_hp_in(2).W.DATA, --[C_SAXIGP4_DATA_WIDTH-1:0]
      saxigp4_wstrb => s_axi_hp_in(2).W.STRB, --[(C_SAXIGP4_DATA_WIDTH/8) -1 :0]
      saxigp4_wlast => s_axi_hp_in(2).W.LAST,
      saxigp4_wvalid => s_axi_hp_in(2).W.VALID,
      saxigp4_wready => s_axi_hp_out(2).W.READY,
      saxigp4_bid => s_axi_hp_out(2).B.ID(5 downto 0), --[5:0]
      saxigp4_bresp => s_axi_hp_out(2).B.RESP, --[1:0]
      saxigp4_bvalid => s_axi_hp_out(2).B.VALID,
      saxigp4_bready => s_axi_hp_in(2).B.READY,
      saxigp4_arid => s_axi_hp_in(2).AR.ID(5 downto 0), --[5:0]
      saxigp4_araddr => saxigp_araddrs(2), --[48:0]
      saxigp4_arlen => saxigp_arlens(2), --[7:0]
      saxigp4_arsize => s_axi_hp_in(2).AR.SIZE, --[2:0]
      saxigp4_arburst => s_axi_hp_in(2).AR.BURST, --[1:0]
      saxigp4_arlock => s_axi_hp_in(2).AR.LOCK(0),
      saxigp4_arcache => s_axi_hp_in(2).AR.CACHE, --[3:0]
      saxigp4_arprot => s_axi_hp_in(2).AR.PROT, --[2:0]
      saxigp4_arvalid => s_axi_hp_in(2).AR.VALID,
      saxigp4_arready => s_axi_hp_out(2).AR.READY,
      saxigp4_rid => s_axi_hp_out(2).R.ID(5 downto 0), --[5:0]
      saxigp4_rdata => s_axi_hp_out(2).R.DATA, --[C_SAXIGP4_DATA_WIDTH-1:0]
      saxigp4_rresp => s_axi_hp_out(2).R.RESP, --[1:0]
      saxigp4_rlast => s_axi_hp_out(2).R.LAST,
      saxigp4_rvalid => s_axi_hp_out(2).R.VALID,
      saxigp4_rready => s_axi_hp_in(2).R.READY,
      saxigp4_awqos => s_axi_hp_in(2).AW.QOS, --[3:0]
      saxigp4_arqos => s_axi_hp_in(2).AR.QOS, --[3:0]
      saxigp4_rcount => s_axi_hp_out(2).R.COUNT, --[7:0]
      saxigp4_wcount => s_axi_hp_out(2).W.COUNT, --[7:0]
      saxigp4_racount => saxigp_racounts(2), --[3:0]
      saxigp4_wacount => s_axi_hp_out(2).AW.COUNT(3 downto 0), --[3:0]
-- saxigp5
      saxihp3_fpd_aclk => s_axi_hp_in(3).ACLK,
      saxihp3_fpd_rclk => '0',
      saxihp3_fpd_wclk => '0',
      saxigp5_aruser => '0',
      saxigp5_awuser => '0',
      saxigp5_awid => s_axi_hp_in(3).AW.ID(5 downto 0), --[5:0]
      saxigp5_awaddr => saxigp_awaddrs(3), --[48:0]
      saxigp5_awlen => saxigp_awlens(3), --[7:0]
      saxigp5_awsize => s_axi_hp_in(3).AW.SIZE, --[2:0]
      saxigp5_awburst => s_axi_hp_in(3).AW.BURST, --[1:0]
      saxigp5_awlock => s_axi_hp_in(3).AW.LOCK(0),
      saxigp5_awcache => s_axi_hp_in(3).AW.CACHE, --[3:0]
      saxigp5_awprot => s_axi_hp_in(3).AW.PROT, --[2:0]
      saxigp5_awvalid => s_axi_hp_in(3).AW.VALID,
      saxigp5_awready => s_axi_hp_out(3).AW.READY,
      saxigp5_wdata => s_axi_hp_in(3).W.DATA, --[C_SAXIGP5_DATA_WIDTH-1:0]
      saxigp5_wstrb => s_axi_hp_in(3).W.STRB, --[(C_SAXIGP5_DATA_WIDTH/8) -1 :0]
      saxigp5_wlast => s_axi_hp_in(3).W.LAST,
      saxigp5_wvalid => s_axi_hp_in(3).W.VALID,
      saxigp5_wready => s_axi_hp_out(3).W.READY,
      saxigp5_bid => s_axi_hp_out(3).B.ID(5 downto 0), --[5:0]
      saxigp5_bresp => s_axi_hp_out(3).B.RESP, --[1:0]
      saxigp5_bvalid => s_axi_hp_out(3).B.VALID,
      saxigp5_bready => s_axi_hp_in(3).B.READY,
      saxigp5_arid => s_axi_hp_in(3).AR.ID(5 downto 0), --[5:0]
      saxigp5_araddr => saxigp_araddrs(3), --[48:0]
      saxigp5_arlen => saxigp_arlens(3), --[7:0]
      saxigp5_arsize => s_axi_hp_in(3).AR.SIZE, --[2:0]
      saxigp5_arburst => s_axi_hp_in(3).AR.BURST, --[1:0]
      saxigp5_arlock => s_axi_hp_in(3).AR.LOCK(0),
      saxigp5_arcache => s_axi_hp_in(3).AR.CACHE, --[3:0]
      saxigp5_arprot => s_axi_hp_in(3).AR.PROT, --[2:0]
      saxigp5_arvalid => s_axi_hp_in(3).AR.VALID,
      saxigp5_arready => s_axi_hp_out(3).AR.READY,
      saxigp5_rid => s_axi_hp_out(3).R.ID(5 downto 0), --[5:0]
      saxigp5_rdata => s_axi_hp_out(3).R.DATA, --[C_SAXIGP5_DATA_WIDTH-1:0]
      saxigp5_rresp => s_axi_hp_out(3).R.RESP, --[1:0]
      saxigp5_rlast => s_axi_hp_out(3).R.LAST,
      saxigp5_rvalid => s_axi_hp_out(3).R.VALID,
      saxigp5_rready => s_axi_hp_in(3).R.READY,
      saxigp5_awqos => s_axi_hp_in(3).AW.QOS, --[3:0]
      saxigp5_arqos => s_axi_hp_in(3).AR.QOS, --[3:0]
      saxigp5_rcount => s_axi_hp_out(3).R.COUNT, --[7:0]
      saxigp5_wcount => s_axi_hp_out(3).W.COUNT, --[7:0]
      saxigp5_racount => saxigp_racounts(3), --[3:0]
      saxigp5_wacount => s_axi_hp_out(3).AW.COUNT(3 downto 0), --[3:0]
-- saxigp6
      --NOT USING
      saxi_lpd_aclk => '0', -- s_axi_hp_in(6).ACLK,
      saxi_lpd_rclk => '0',
      saxi_lpd_wclk => '0',
      saxigp6_aruser => '0', -- s_axi_hp_in(6).ARUSER,
      saxigp6_awuser => '0', -- s_axi_hp_in(6).AWUSER,
      saxigp6_awid => (others => '0'), -- s_axi_hp_in(6).AW.ID, --[5:0]
      saxigp6_awaddr => (others => '0'), -- s_axi_hp_in(6).AW.ADDR, --[48:0]
      saxigp6_awlen => (others => '0'), -- s_axi_hp_in(6).AW.LEN, --[7:0]
      saxigp6_awsize => (others => '0'), -- s_axi_hp_in(6).AW.SIZE, --[2:0]
      saxigp6_awburst => (others => '0'), -- s_axi_hp_in(6).AW.BURST, --[1:0]
      saxigp6_awlock => '0', -- s_axi_hp_in(6).AW.LOCK(0),
      saxigp6_awcache => (others => '0'), -- s_axi_hp_in(6).AW.CACHE, --[3:0]
      saxigp6_awprot => (others => '0'), -- s_axi_hp_in(6).AW.PROT, --[2:0]
      saxigp6_awvalid => '0', -- s_axi_hp_in(6).AW.VALID,
      saxigp6_awready => open, -- s_axi_hp_out(6).AW.READY,
      saxigp6_wdata => (others => '0'), -- s_axi_hp_in(6).W.DATA, --[C_SAXIGP6_DATA_WIDTH-1:0]
      saxigp6_wstrb => (others => '0'), -- s_axi_hp_in(6).W.STRB, --[(C_SAXIGP6_DATA_WIDTH/8) -1 :0]
      saxigp6_wlast => '0', -- s_axi_hp_in(6).W.LAST,
      saxigp6_wvalid => '0', -- s_axi_hp_in(6).W.VALID,
      saxigp6_wready => open, -- s_axi_hp_out(6).W.READY,
      saxigp6_bid => open, -- s_axi_hp_out(6).B.ID, --[5:0]
      saxigp6_bresp => open, -- s_axi_hp_out(6).B.RESP, --[1:0]
      saxigp6_bvalid => open, -- s_axi_hp_out(6).B.VALID,
      saxigp6_bready => '0', -- s_axi_hp_in(6).B.READY,
      saxigp6_arid => (others => '0'), -- s_axi_hp_in(6).AR.ID, --[5:0]
      saxigp6_araddr => (others => '0'), -- s_axi_hp_in(6).AR.ADDR, --[48:0]
      saxigp6_arlen => (others => '0'), -- s_axi_hp_in(6).AR.LEN, --[7:0]
      saxigp6_arsize => (others => '0'), -- s_axi_hp_in(6).AR.SIZE, --[2:0]
      saxigp6_arburst => (others => '0'), -- s_axi_hp_in(6).AR.BURST, --[1:0]
      saxigp6_arlock => '0', -- s_axi_hp_in(6).AR.LOCK(0),
      saxigp6_arcache => (others => '0'), -- s_axi_hp_in(6).AR.CACHE, --[3:0]
      saxigp6_arprot => (others => '0'), -- s_axi_hp_in(6).AR.PROT, --[2:0]
      saxigp6_arvalid => '0', -- s_axi_hp_in(6).AR.VALID,
      saxigp6_arready => open, -- s_axi_hp_out(6).AR.READY,
      saxigp6_rid => open, -- s_axi_hp_out(6).R.ID, --[5:0]
      saxigp6_rdata => open, -- s_axi_hp_out(6).R.DATA, --[C_SAXIGP6_DATA_WIDTH-1:0]
      saxigp6_rresp => open, -- s_axi_hp_out(6).R.RESP, --[1:0]
      saxigp6_rlast => open, -- s_axi_hp_out(6).R.LAST,
      saxigp6_rvalid => open, -- s_axi_hp_out(6).R.VALID,
      saxigp6_rready => '0', -- s_axi_hp_in(6).R.READY,
      saxigp6_awqos => (others => '0'), -- s_axi_hp_in(6).AW.QOS, --[3:0]
      saxigp6_arqos => (others => '0'), -- s_axi_hp_in(6).AR.QOS, --[3:0]
      saxigp6_rcount => open, -- s_axi_hp_out(6).R.COUNT, --[7:0]
      saxigp6_wcount => open, -- s_axi_hp_out(6).W.COUNT, --[7:0]
      saxigp6_racount => open, -- s_axi_hp_out(6).AR.COUNT, --[3:0]
      saxigp6_wacount => open, -- s_axi_hp_out(6).AW.COUNT, --[3:0]
-- saxiacp
      -- NOT USING
      saxiacp_fpd_aclk => '0',
      saxiacp_awaddr => (others => '0'), --[39:0]
      saxiacp_awid => (others => '0'), --[4:0]
      saxiacp_awlen => (others => '0'), --[7:0]
      saxiacp_awsize => (others => '0'), --[2:0]
      saxiacp_awburst => (others => '0'), --[1:0]
      saxiacp_awlock => '0',
      saxiacp_awcache => (others => '0'), --[3:0]
      saxiacp_awprot => (others => '0'), --[2:0]
      saxiacp_awvalid => '0',
      saxiacp_awready => open,
      saxiacp_awuser => (others => '0'), --[1:0]
      saxiacp_awqos => (others => '0'), --[3:0]
      saxiacp_wlast => '0',
      saxiacp_wdata => (others => '0'), --[127:0]
      saxiacp_wstrb => (others => '0'), --[15:0]
      saxiacp_wvalid => '0',
      saxiacp_wready => open,
      saxiacp_bresp => open, --[1:0]
      saxiacp_bid => open, --[4:0]
      saxiacp_bvalid => open,
      saxiacp_bready => '0',
      saxiacp_araddr => (others => '0'), --[39:0]
      saxiacp_arid => (others => '0'), --[4:0]
      saxiacp_arlen => (others => '0'), --[7:0]
      saxiacp_arsize => (others => '0'), --[2:0]
      saxiacp_arburst => (others => '0'), --[1:0]
      saxiacp_arlock => '0',
      saxiacp_arcache => (others => '0'), --[3:0]
      saxiacp_arprot => (others => '0'), --[2:0]
      saxiacp_arvalid => '0',
      saxiacp_arready => open,
      saxiacp_aruser => (others => '0'), --[1:0]
      saxiacp_arqos => (others => '0'), --[3:0]
      saxiacp_rid => open, --[4:0]
      saxiacp_rlast => open,
      saxiacp_rdata => open, --[127:0]
      saxiacp_rresp => open, --[1:0]
      saxiacp_rvalid => open,
      saxiacp_rready => '0',
-- sacefpd
      -- NOT USING
      sacefpd_aclk => '0',
      sacefpd_awvalid => '0',
      sacefpd_awready => open,
      sacefpd_awid => (others => '0'), --[5:0]
      sacefpd_awaddr => (others => '0'), --[43:0]
      sacefpd_awregion => (others => '0'), --[3:0]
      sacefpd_awlen => (others => '0'), --[7:0]
      sacefpd_awsize => (others => '0'), --[2:0]
      sacefpd_awburst => (others => '0'), --[1:0]
      sacefpd_awlock => '0',
      sacefpd_awcache => (others => '0'), --[3:0]
      sacefpd_awprot => (others => '0'), --[2:0]
      sacefpd_awdomain => (others => '0'), --[1:0]
      sacefpd_awsnoop => (others => '0'), --[2:0]
      sacefpd_awbar => (others => '0'), --[1:0]
      sacefpd_awqos => (others => '0'), --[3:0]
      sacefpd_wvalid => '0',
      sacefpd_wready => open,
      sacefpd_wdata => (others => '0'), --[127:0]
      sacefpd_wstrb => (others => '0'), --[15:0]
      sacefpd_wlast => '0',
      sacefpd_wuser => '0',
      sacefpd_bvalid => open,
      sacefpd_bready => '0',
      sacefpd_bid => open, --[5:0]
      sacefpd_bresp => open, --[1:0]
      sacefpd_buser => open,
      sacefpd_arvalid => '0',
      sacefpd_arready => open,
      sacefpd_arid => (others => '0'), --[5:0]
      sacefpd_araddr => (others => '0'), --[43:0]
      sacefpd_arregion => (others => '0'), --[3:0]
      sacefpd_arlen => (others => '0'), --[7:0]
      sacefpd_arsize => (others => '0'), --[2:0]
      sacefpd_arburst => (others => '0'), --[1:0]
      sacefpd_arlock => '0',
      sacefpd_arcache => (others => '0'), --[3:0]
      sacefpd_arprot => (others => '0'), --[2:0]
      sacefpd_ardomain => (others => '0'), --[1:0]
      sacefpd_arsnoop => (others => '0'), --[3:0]
      sacefpd_arbar => (others => '0'), --[1:0]
      sacefpd_arqos => (others => '0'), --[3:0]
      sacefpd_rvalid => open,
      sacefpd_rready => '0',
      sacefpd_rid => open, --[5:0]
      sacefpd_rdata => open, --[127:0]
      sacefpd_rresp => open, --[3:0]
      sacefpd_rlast => open,
      sacefpd_ruser => open,
      sacefpd_acvalid => open,
      sacefpd_acready => '0',
      sacefpd_acaddr => open, --[43:0]
      sacefpd_acsnoop => open, --[3:0]
      sacefpd_acprot => open, --[2:0]
      sacefpd_crvalid => '0',
      sacefpd_crready => open,
      sacefpd_crresp => (others => '0'), --[4:0]
      sacefpd_cdvalid => '0',
      sacefpd_cdready => open,
      sacefpd_cddata => (others => '0'), --[127:0]
      sacefpd_cdlast => '0',
      sacefpd_wack => '0',
      sacefpd_rack => '0',


-----------------------------------------------
-- not using anything below this line yet... --
-----------------------------------------------

-- can0
      emio_can0_phy_tx => open,
      emio_can0_phy_rx => '0',
-- can1
      emio_can1_phy_tx => open,
      emio_can1_phy_rx => '0',
-- enet0
      emio_enet0_gmii_rx_clk => '0',
      emio_enet0_speed_mode => open, --[2:0]
      emio_enet0_gmii_crs => '0',
      emio_enet0_gmii_col => '0',
      emio_enet0_gmii_rxd => (others => '0'), --[7:0]
      emio_enet0_gmii_rx_er => '0',
      emio_enet0_gmii_rx_dv => '0',
      emio_enet0_gmii_tx_clk => '0',
      emio_enet0_gmii_txd => open, --[7:0]
      emio_enet0_gmii_tx_en => open,
      emio_enet0_gmii_tx_er => open,
      emio_enet0_mdio_mdc => open,
      emio_enet0_mdio_i => '0',
      emio_enet0_mdio_o => open,
      emio_enet0_mdio_t => open,
      emio_enet0_mdio_t_n => open,
-- enet1
      emio_enet1_gmii_rx_clk => '0',
      emio_enet1_speed_mode => open, --[2:0]
      emio_enet1_gmii_crs => '0',
      emio_enet1_gmii_col => '0',
      emio_enet1_gmii_rxd => (others => '0'), --[7:0]
      emio_enet1_gmii_rx_er => '0',
      emio_enet1_gmii_rx_dv => '0',
      emio_enet1_gmii_tx_clk => '0',
      emio_enet1_gmii_txd => open, --[7:0]
      emio_enet1_gmii_tx_en => open,
      emio_enet1_gmii_tx_er => open,
      emio_enet1_mdio_mdc => open,
      emio_enet1_mdio_i => '0',
      emio_enet1_mdio_o => open,
      emio_enet1_mdio_t => open,
      emio_enet1_mdio_t_n => open,
-- enet2
      emio_enet2_gmii_rx_clk => '0',
      emio_enet2_speed_mode => open, --[2:0]
      emio_enet2_gmii_crs => '0',
      emio_enet2_gmii_col => '0',
      emio_enet2_gmii_rxd => (others => '0'), --[7:0]
      emio_enet2_gmii_rx_er => '0',
      emio_enet2_gmii_rx_dv => '0',
      emio_enet2_gmii_tx_clk => '0',
      emio_enet2_gmii_txd => open, --[7:0]
      emio_enet2_gmii_tx_en => open,
      emio_enet2_gmii_tx_er => open,
      emio_enet2_mdio_mdc => open,
      emio_enet2_mdio_i => '0',
      emio_enet2_mdio_o => open,
      emio_enet2_mdio_t => open,
      emio_enet2_mdio_t_n => open,
-- enet3
      emio_enet3_gmii_rx_clk => '0',
      emio_enet3_speed_mode => open, --[2:0]
      emio_enet3_gmii_crs => '0',
      emio_enet3_gmii_col => '0',
      emio_enet3_gmii_rxd => (others => '0'), --[7:0]
      emio_enet3_gmii_rx_er => '0',
      emio_enet3_gmii_rx_dv => '0',
      emio_enet3_gmii_tx_clk => '0',
      emio_enet3_gmii_txd => open, --[7:0]
      emio_enet3_gmii_tx_en => open,
      emio_enet3_gmii_tx_er => open,
      emio_enet3_mdio_mdc => open,
      emio_enet3_mdio_i => '0',
      emio_enet3_mdio_o => open,
      emio_enet3_mdio_t => open,
      emio_enet3_mdio_t_n => open,
-- fifoif0
      emio_enet0_tx_r_data_rdy => '0',
      emio_enet0_tx_r_rd => open,
      emio_enet0_tx_r_valid => '0',
      emio_enet0_tx_r_data => (others => '0'), --[7:0]
      emio_enet0_tx_r_sop => '0',
      emio_enet0_tx_r_eop => '0',
      emio_enet0_tx_r_err => '0',
      emio_enet0_tx_r_underflow => '0',
      emio_enet0_tx_r_flushed => '0',
      emio_enet0_tx_r_control => '0',
      emio_enet0_dma_tx_end_tog => open,
      emio_enet0_dma_tx_status_tog => '0',
      emio_enet0_tx_r_status => open, --[3:0]
      emio_enet0_rx_w_wr => open,
      emio_enet0_rx_w_data => open, --[7:0]
      emio_enet0_rx_w_sop => open,
      emio_enet0_rx_w_eop => open,
      emio_enet0_rx_w_status => open, --[44:0]
      emio_enet0_rx_w_err => open,
      emio_enet0_rx_w_overflow => '0',
      emio_enet0_signal_detect => '0',
      emio_enet0_rx_w_flush => open,
      emio_enet0_tx_r_fixed_lat => open,
-- fifoif1
      emio_enet1_tx_r_data_rdy => '0',
      emio_enet1_tx_r_rd => open,
      emio_enet1_tx_r_valid => '0',
      emio_enet1_tx_r_data => (others => '0'), --[7:0]
      emio_enet1_tx_r_sop => '0',
      emio_enet1_tx_r_eop => '0',
      emio_enet1_tx_r_err => '0',
      emio_enet1_tx_r_underflow => '0',
      emio_enet1_tx_r_flushed => '0',
      emio_enet1_tx_r_control => '0',
      emio_enet1_dma_tx_end_tog => open,
      emio_enet1_dma_tx_status_tog => '0',
      emio_enet1_tx_r_status => open, --[3:0]
      emio_enet1_rx_w_wr => open,
      emio_enet1_rx_w_data => open, --[7:0]
      emio_enet1_rx_w_sop => open,
      emio_enet1_rx_w_eop => open,
      emio_enet1_rx_w_status => open, --[44:0]
      emio_enet1_rx_w_err => open,
      emio_enet1_rx_w_overflow => '0',
      emio_enet1_signal_detect => '0',
      emio_enet1_rx_w_flush => open,
      emio_enet1_tx_r_fixed_lat => open,
-- fifoif2
      emio_enet2_tx_r_data_rdy => '0',
      emio_enet2_tx_r_rd => open,
      emio_enet2_tx_r_valid => '0',
      emio_enet2_tx_r_data => (others => '0'), --[7:0]
      emio_enet2_tx_r_sop => '0',
      emio_enet2_tx_r_eop => '0',
      emio_enet2_tx_r_err => '0',
      emio_enet2_tx_r_underflow => '0',
      emio_enet2_tx_r_flushed => '0',
      emio_enet2_tx_r_control => '0',
      emio_enet2_dma_tx_end_tog => open,
      emio_enet2_dma_tx_status_tog => '0',
      emio_enet2_tx_r_status => open, --[3:0]
      emio_enet2_rx_w_wr => open,
      emio_enet2_rx_w_data => open, --[7:0]
      emio_enet2_rx_w_sop => open,
      emio_enet2_rx_w_eop => open,
      emio_enet2_rx_w_status => open, --[44:0]
      emio_enet2_rx_w_err => open,
      emio_enet2_rx_w_overflow => '0',
      emio_enet2_signal_detect => '0',
      emio_enet2_rx_w_flush => open,
      emio_enet2_tx_r_fixed_lat => open,
-- fifoif3
      emio_enet3_tx_r_data_rdy => '0',
      emio_enet3_tx_r_rd => open,
      emio_enet3_tx_r_valid => '0',
      emio_enet3_tx_r_data => (others => '0'), --[7:0]
      emio_enet3_tx_r_sop => '0',
      emio_enet3_tx_r_eop => '0',
      emio_enet3_tx_r_err => '0',
      emio_enet3_tx_r_underflow => '0',
      emio_enet3_tx_r_flushed => '0',
      emio_enet3_tx_r_control => '0',
      emio_enet3_dma_tx_end_tog => open,
      emio_enet3_dma_tx_status_tog => '0',
      emio_enet3_tx_r_status => open, --[3:0]
      emio_enet3_rx_w_wr => open,
      emio_enet3_rx_w_data => open, --[7:0]
      emio_enet3_rx_w_sop => open,
      emio_enet3_rx_w_eop => open,
      emio_enet3_rx_w_status => open, --[44:0]
      emio_enet3_rx_w_err => open,
      emio_enet3_rx_w_overflow => '0',
      emio_enet3_signal_detect => '0',
      emio_enet3_rx_w_flush => open,
      emio_enet3_tx_r_fixed_lat => open,
-- gem0_fmio
--      fmio_gem0_fifo_tx_clk_from_pl => '0',
--      fmio_gem0_fifo_rx_clk_from_pl => '0',
      fmio_gem0_fifo_tx_clk_to_pl_bufg => open,
      fmio_gem0_fifo_rx_clk_to_pl_bufg => open,
-- gem1_fmio
--      fmio_gem1_fifo_tx_clk_from_pl => '0',
--      fmio_gem1_fifo_rx_clk_from_pl => '0',
      fmio_gem1_fifo_tx_clk_to_pl_bufg => open,
      fmio_gem1_fifo_rx_clk_to_pl_bufg => open,
-- gem2_fmio
--      fmio_gem2_fifo_tx_clk_from_pl => '0',
--      fmio_gem2_fifo_rx_clk_from_pl => '0',
      fmio_gem2_fifo_tx_clk_to_pl_bufg => open,
      fmio_gem2_fifo_rx_clk_to_pl_bufg => open,
-- gem3_fmio
--      fmio_gem3_fifo_tx_clk_from_pl => '0',
--      fmio_gem3_fifo_rx_clk_from_pl => '0',
      fmio_gem3_fifo_tx_clk_to_pl_bufg => open,
      fmio_gem3_fifo_rx_clk_to_pl_bufg => open,
-- gem0_1588
       emio_enet0_tx_sof => open,
       emio_enet0_sync_frame_tx => open,
       emio_enet0_delay_req_tx => open,
       emio_enet0_pdelay_req_tx => open,
       emio_enet0_pdelay_resp_tx => open,
       emio_enet0_rx_sof => open,
       emio_enet0_sync_frame_rx => open,
       emio_enet0_delay_req_rx => open,
       emio_enet0_pdelay_req_rx => open,
       emio_enet0_pdelay_resp_rx => open,
       emio_enet0_tsu_inc_ctrl => (others => '0'), --[1:0]
       emio_enet0_tsu_timer_cmp_val => open,
--gem1_1588
       emio_enet1_tx_sof => open,
       emio_enet1_sync_frame_tx => open,
       emio_enet1_delay_req_tx => open,
       emio_enet1_pdelay_req_tx => open,
       emio_enet1_pdelay_resp_tx => open,
       emio_enet1_rx_sof => open,
       emio_enet1_sync_frame_rx => open,
       emio_enet1_delay_req_rx => open,
       emio_enet1_pdelay_req_rx => open,
       emio_enet1_pdelay_resp_rx => open,
       emio_enet1_tsu_inc_ctrl => (others => '0'), --[1:0]
       emio_enet1_tsu_timer_cmp_val => open,
--gem2_1588
       emio_enet2_tx_sof => open,
       emio_enet2_sync_frame_tx => open,
       emio_enet2_delay_req_tx => open,
       emio_enet2_pdelay_req_tx => open,
       emio_enet2_pdelay_resp_tx => open,
       emio_enet2_rx_sof => open,
       emio_enet2_sync_frame_rx => open,
       emio_enet2_delay_req_rx => open,
       emio_enet2_pdelay_req_rx => open,
       emio_enet2_pdelay_resp_rx => open,
       emio_enet2_tsu_inc_ctrl => (others => '0'), --[1:0]
       emio_enet2_tsu_timer_cmp_val => open,
--gem3_1588
       emio_enet3_tx_sof => open,
       emio_enet3_sync_frame_tx => open,
       emio_enet3_delay_req_tx => open,
       emio_enet3_pdelay_req_tx => open,
       emio_enet3_pdelay_resp_tx => open,
       emio_enet3_rx_sof => open,
       emio_enet3_sync_frame_rx => open,
       emio_enet3_delay_req_rx => open,
       emio_enet3_pdelay_req_rx => open,
       emio_enet3_pdelay_resp_rx => open,
       emio_enet3_tsu_inc_ctrl => (others => '0'), --[1:0]
       emio_enet3_tsu_timer_cmp_val => open,
-- gem_tsu
      fmio_gem_tsu_clk_from_pl => '0',
      fmio_gem_tsu_clk_to_pl_bufg => open,
      emio_enet_tsu_clk => '0',
      emio_enet0_enet_tsu_timer_cnt => open, --[93:0]
-- gem_misc
      emio_enet0_ext_int_in => '0',
      emio_enet1_ext_int_in => '0',
      emio_enet2_ext_int_in => '0',
      emio_enet3_ext_int_in => '0',
      emio_enet0_dma_bus_width => open, --[1:0]
      emio_enet1_dma_bus_width => open, --[1:0]
      emio_enet2_dma_bus_width => open, --[1:0]
      emio_enet3_dma_bus_width => open, --[1:0]
-- gpio
      emio_gpio_i => (others => '0'), --[(C_EMIO_GPIO_WIDTH -1):0]
      emio_gpio_o => open, --[(C_EMIO_GPIO_WIDTH -1):0]
      emio_gpio_t => open, --[(C_EMIO_GPIO_WIDTH -1):0]
      emio_gpio_t_n => open, --[(C_EMIO_GPIO_WIDTH -1):0]
-- i2c0
      emio_i2c0_scl_i => '0',
      emio_i2c0_scl_o => open,
      emio_i2c0_scl_t_n => open,
      emio_i2c0_scl_t => open,
      emio_i2c0_sda_i => '0',
      emio_i2c0_sda_o => open,
      emio_i2c0_sda_t_n => open,
      emio_i2c0_sda_t => open,
-- i2c1
      emio_i2c1_scl_i => '0',
      emio_i2c1_scl_o => open,
      emio_i2c1_scl_t => open,
      emio_i2c1_scl_t_n => open,
      emio_i2c1_sda_i => '0',
      emio_i2c1_sda_o => open,
      emio_i2c1_sda_t => open,
      emio_i2c1_sda_t_n => open,
-- uart0
      emio_uart0_txd => open,
      emio_uart0_rxd => '0',
      emio_uart0_ctsn => '0',
      emio_uart0_rtsn => open,
      emio_uart0_dsrn => '0',
      emio_uart0_dcdn => '0',
      emio_uart0_rin => '0',
      emio_uart0_dtrn => open,
-- uart1
      emio_uart1_txd => open,
      emio_uart1_rxd => '0',
      emio_uart1_ctsn => '0',
      emio_uart1_rtsn => open,
      emio_uart1_dsrn => '0',
      emio_uart1_dcdn => '0',
      emio_uart1_rin => '0',
      emio_uart1_dtrn => open,
-- sdio0
      emio_sdio0_clkout => open,
      emio_sdio0_fb_clk_in => '0',
      emio_sdio0_cmdout => open,
      emio_sdio0_cmdin => '0',
      emio_sdio0_cmdena => open,
      emio_sdio0_datain => (others => '0'), --[C_SD0_INTERNAL_BUS_WIDTH-1:0]
      emio_sdio0_dataout => open, --[C_SD0_INTERNAL_BUS_WIDTH-1:0]
      emio_sdio0_dataena => open, --[C_SD0_INTERNAL_BUS_WIDTH-1:0]
      emio_sdio0_cd_n => '0',
      emio_sdio0_wp => '0',
      emio_sdio0_ledcontrol => open,
      emio_sdio0_buspower => open,
      emio_sdio0_bus_volt => open, --[2:0]
-- sdio1
      emio_sdio1_clkout => open,
      emio_sdio1_fb_clk_in => '0',
      emio_sdio1_cmdout => open,
      emio_sdio1_cmdin => '0',
      emio_sdio1_cmdena => open,
      emio_sdio1_datain => (others => '0'), --[C_SD1_INTERNAL_BUS_WIDTH-1:0]
      emio_sdio1_dataout => open, --[C_SD1_INTERNAL_BUS_WIDTH-1:0]
      emio_sdio1_dataena => open, --[C_SD1_INTERNAL_BUS_WIDTH-1:0]
      emio_sdio1_cd_n => '0',
      emio_sdio1_wp => '0',
      emio_sdio1_ledcontrol => open,
      emio_sdio1_buspower => open,
      emio_sdio1_bus_volt => open, --[2:0]
-- spi0
      emio_spi0_sclk_i => '0',
      emio_spi0_sclk_o => open,
      emio_spi0_sclk_t => open,
      emio_spi0_sclk_t_n => open,
      emio_spi0_m_i => '0',
      emio_spi0_m_o => open,
      emio_spi0_mo_t => open,
      emio_spi0_mo_t_n => open,
      emio_spi0_s_i => '0',
      emio_spi0_s_o => open,
      emio_spi0_so_t => open,
      emio_spi0_so_t_n => open,
      emio_spi0_ss_i_n => '0',
      emio_spi0_ss_o_n => open,
      emio_spi0_ss1_o_n => open,
      emio_spi0_ss2_o_n => open,
      emio_spi0_ss_n_t => open,
      emio_spi0_ss_n_t_n => open,
-- spi1
      emio_spi1_sclk_i => '0',
      emio_spi1_sclk_o => open,
      emio_spi1_sclk_t => open,
      emio_spi1_sclk_t_n => open,
      emio_spi1_m_i => '0',
      emio_spi1_m_o => open,
      emio_spi1_mo_t => open,
      emio_spi1_mo_t_n => open,
      emio_spi1_s_i => '0',
      emio_spi1_s_o => open,
      emio_spi1_so_t => open,
      emio_spi1_so_t_n => open,
      emio_spi1_ss_i_n => '0',
      emio_spi1_ss_o_n => open,
      emio_spi1_ss1_o_n => open,
      emio_spi1_ss2_o_n => open,
      emio_spi1_ss_n_t => open,
      emio_spi1_ss_n_t_n => open,
-- trace
      pl_ps_trace_clk => '0',
      ps_pl_tracectl => open,
      ps_pl_tracedata => open, --[C_TRACE_DATA_WIDTH-1:0]
      trace_clk_out => open,
-- ttc0
      emio_ttc0_wave_o => open, --[2:0]
      emio_ttc0_clk_i => (others => '0'), --[2:0]
-- ttc1
      emio_ttc1_wave_o => open, --[2:0]
      emio_ttc1_clk_i => (others => '0'), --[2:0]
-- ttc2
      emio_ttc2_wave_o => open, --[2:0]
      emio_ttc2_clk_i => (others => '0'), --[2:0]
-- ttc3
      emio_ttc3_wave_o => open, --[2:0]
      emio_ttc3_clk_i => (others => '0'), --[2:0]
-- wdt0
      emio_wdt0_clk_i => '0',
      emio_wdt0_rst_o => open,
-- wdt1
      emio_wdt1_clk_i => '0',
      emio_wdt1_rst_o => open,
-- usb3
      emio_hub_port_overcrnt_usb3_0 => '0',
      emio_hub_port_overcrnt_usb3_1 => '0',
      emio_hub_port_overcrnt_usb2_0 => '0',
      emio_hub_port_overcrnt_usb2_1 => '0',
      emio_u2dsport_vbus_ctrl_usb3_0 => open,
      emio_u2dsport_vbus_ctrl_usb3_1 => open,
      emio_u3dsport_vbus_ctrl_usb3_0 => open,
      emio_u3dsport_vbus_ctrl_usb3_1 => open,
--adma
      adma_fci_clk => (others => '0'), --[7:0]
      pl2adma_cvld => (others => '0'), --[7:0]
      pl2adma_tack => (others => '0'), --[7:0]
      adma2pl_cack => open, --[7:0]
      adma2pl_tvld => open, --[7:0]
--gdma
      perif_gdma_clk => (others => '0'), --[7:0]
      perif_gdma_cvld => (others => '0'), --[7:0]
      perif_gdma_tack => (others => '0'), --[7:0]
      gdma_perif_cack => open, --[7:0]
      gdma_perif_tvld => open, --[7:0]
-- clk
      pl_clock_stop => (others => '0'), --[3:0]
      pll_aux_refclk_lpd => (others => '0'), --[1:0]
      pll_aux_refclk_fpd => (others => '0'), --[2:0]
-- audio
      dp_s_axis_audio_tdata => (others => '0'), --[31:0]
      dp_s_axis_audio_tid => '0',
      dp_s_axis_audio_tvalid => '0',
      dp_s_axis_audio_tready => open,
      dp_m_axis_mixed_audio_tdata => open, --[31:0]
      dp_m_axis_mixed_audio_tid => open,
      dp_m_axis_mixed_audio_tvalid => open,
      dp_m_axis_mixed_audio_tready => '0',
      dp_s_axis_audio_clk => '0',
-- video
      dp_live_video_in_vsync => '0',
      dp_live_video_in_hsync => '0',
      dp_live_video_in_de => '0',
      dp_live_video_in_pixel1 => (others => '0'), --[35:0]
      dp_video_in_clk => '0',
      dp_video_out_hsync => open,
      dp_video_out_vsync => open,
      dp_video_out_pixel1 => open, --[35:0]
      dp_aux_data_in => '0',
      dp_aux_data_out => open,
      dp_aux_data_oe_n => open,
      dp_live_gfx_alpha_in => (others => '0'), --[7:0]
      dp_live_gfx_pixel1_in => (others => '0'), --[35:0]
      dp_hot_plug_detect => '0',
      dp_external_custom_event1 => '0',
      dp_external_custom_event2 => '0',
      dp_external_vsync_event => '0',
      dp_live_video_de_out => open,
-- event_apu
      pl_ps_eventi => '0',
      ps_pl_evento => open,
      ps_pl_standbywfe => open, --[3:0]
      ps_pl_standbywfi => open, --[3:0]
      pl_ps_apugic_irq => (others => '0'), --[3:0]
      pl_ps_apugic_fiq => (others => '0'), --[3:0]
-- event_rpu
      rpu_eventi0 => '0',
      rpu_eventi1 => '0',
      rpu_evento0 => open,
      rpu_evento1 => open,
      nfiq0_lpd_rpu => '0',
      nfiq1_lpd_rpu => '0',
      nirq0_lpd_rpu => '0',
      nirq1_lpd_rpu => '0',
-- ipi
      irq_ipi_pl_0 => open,
      irq_ipi_pl_1 => open,
      irq_ipi_pl_2 => open,
      irq_ipi_pl_3 => open,
-- stm
      stm_event => (others => '0'), --[59:0]
-- ftm
      pl_ps_trigack_0 => '0',
      pl_ps_trigack_1 => '0',
      pl_ps_trigack_2 => '0',
      pl_ps_trigack_3 => '0',
      pl_ps_trigger_0 => '0',
      pl_ps_trigger_1 => '0',
      pl_ps_trigger_2 => '0',
      pl_ps_trigger_3 => '0',
      ps_pl_trigack_0 => open,
      ps_pl_trigack_1 => open,
      ps_pl_trigack_2 => open,
      ps_pl_trigack_3 => open,
      ps_pl_trigger_0 => open,
      ps_pl_trigger_1 => open,
      ps_pl_trigger_2 => open,
      ps_pl_trigger_3 => open,
      ftm_gpo => open, --[31:0]
      ftm_gpi => ps_in.debug, -- (others => '0'), --[31:0]
-- irq
      pl_ps_irq0 => (others => '0'), --[(C_NUM_F2P_0_INTR_INPUTS-1):0]
      pl_ps_irq1 => (others => '0'), --[(C_NUM_F2P_1_INTR_INPUTS-1):0]
--      ps_pl_irq_lpd => open, --[99:0]
--      ps_pl_irq_fpd => open, --[63:0]

--resets using gpio

      pl_resetn0 => ps_out.FCLKRESET_N,
      pl_resetn1 => open,
      pl_resetn2 => open,
      pl_resetn3 => open,

      ps_pl_irq_can0 => open,
      ps_pl_irq_can1 => open,
      ps_pl_irq_enet0 => open,
      ps_pl_irq_enet1 => open,
      ps_pl_irq_enet2 => open,
      ps_pl_irq_enet3 => open,
      ps_pl_irq_enet0_wake => open,
      ps_pl_irq_enet1_wake => open,
      ps_pl_irq_enet2_wake => open,
      ps_pl_irq_enet3_wake => open,
      ps_pl_irq_gpio => open,
      ps_pl_irq_i2c0 => open,
      ps_pl_irq_i2c1 => open,
      ps_pl_irq_uart0 => open,
      ps_pl_irq_uart1 => open,
      ps_pl_irq_sdio0 => open,
      ps_pl_irq_sdio1 => open,
      ps_pl_irq_sdio0_wake => open,
      ps_pl_irq_sdio1_wake => open,
      ps_pl_irq_spi0 => open,
      ps_pl_irq_spi1 => open,
      ps_pl_irq_qspi => open,
      ps_pl_irq_ttc0_0 => open,
      ps_pl_irq_ttc0_1 => open,
      ps_pl_irq_ttc0_2 => open,
      ps_pl_irq_ttc1_0 => open,
      ps_pl_irq_ttc1_1 => open,
      ps_pl_irq_ttc1_2 => open,
      ps_pl_irq_ttc2_0 => open,
      ps_pl_irq_ttc2_1 => open,
      ps_pl_irq_ttc2_2 => open,
      ps_pl_irq_ttc3_0 => open,
      ps_pl_irq_ttc3_1 => open,
      ps_pl_irq_ttc3_2 => open,
      ps_pl_irq_csu_pmu_wdt => open,
      ps_pl_irq_lp_wdt => open,
      ps_pl_irq_usb3_0_endpoint => open, --[3:0]
      ps_pl_irq_usb3_0_otg => open,
      ps_pl_irq_usb3_1_endpoint => open, --[3:0]
      ps_pl_irq_usb3_1_otg => open,
      ps_pl_irq_adma_chan => open, --[7:0]
      ps_pl_irq_usb3_0_pmu_wakeup => open, --[1:0]
      ps_pl_irq_gdma_chan => open, --[7:0]
      ps_pl_irq_csu => open,
      ps_pl_irq_csu_dma => open,
      ps_pl_irq_efuse => open,
      ps_pl_irq_xmpu_lpd => open,
      ps_pl_irq_ddr_ss => open,
      ps_pl_irq_nand => open,
      ps_pl_irq_fp_wdt => open,
      ps_pl_irq_pcie_msi => open, --[1:0]
      ps_pl_irq_pcie_legacy => open,
      ps_pl_irq_pcie_dma => open,
      ps_pl_irq_pcie_msc => open,
      ps_pl_irq_dport => open,
      ps_pl_irq_fpd_apb_int => open,
      ps_pl_irq_fpd_atb_error => open,
      ps_pl_irq_dpdma => open,
      ps_pl_irq_apm_fpd => open,
      ps_pl_irq_gpu => open,
      ps_pl_irq_sata => open,
      ps_pl_irq_xmpu_fpd => open,
      ps_pl_irq_apu_cpumnt => open, --[3:0]
      ps_pl_irq_apu_cti => open, --[3:0]
      ps_pl_irq_apu_pmu => open, --[3:0]
      ps_pl_irq_apu_comm => open, --[3:0]
      ps_pl_irq_apu_l2err => open,
      ps_pl_irq_apu_exterr => open,
      ps_pl_irq_apu_regs => open,
      ps_pl_irq_intf_ppd_cci => open,
      ps_pl_irq_intf_fpd_smmu => open,
      ps_pl_irq_atb_err_lpd => open,
      ps_pl_irq_aib_axi => open,
      ps_pl_irq_ams => open,
      ps_pl_irq_lpd_apm => open,
      ps_pl_irq_rtc_alaram => open,
      ps_pl_irq_rtc_seconds => open,
      ps_pl_irq_clkmon => open,
      ps_pl_irq_ipi_channel0 => open,
      ps_pl_irq_ipi_channel1 => open,
      ps_pl_irq_ipi_channel2 => open,
      ps_pl_irq_ipi_channel7 => open,
      ps_pl_irq_ipi_channel8 => open,
      ps_pl_irq_ipi_channel9 => open,
      ps_pl_irq_ipi_channel10 => open,
      ps_pl_irq_rpu_pm => open, --[1:0]
      ps_pl_irq_ocm_error => open,
      ps_pl_irq_lpd_apb_intr => open,
      ps_pl_irq_r5_core0_ecc_error => open,
      ps_pl_irq_r5_core1_ecc_error => open,


-- rtc
      osc_rtc_clk => open,
-- pmu
      pl_pmu_gpi => (others => '0'), --[31:0]
      pmu_pl_gpo => open, --[31:0]
      aib_pmu_afifm_fpd_ack => '0',
      aib_pmu_afifm_lpd_ack => '0',
      pmu_aib_afifm_fpd_req => open,
      pmu_aib_afifm_lpd_req => open,
      pmu_error_to_pl => open, --[46:0]
      pmu_error_from_pl => (others => '0'), --[3:0]
-- misc
      ddrc_ext_refresh_rank0_req => '0',
      ddrc_ext_refresh_rank1_req => '0',
      ddrc_refresh_pl_clk => '0',
      pl_acpinact => '0',

--For Clock buffering
--FCLK
      pl_clk3 => ps_out.FCLK(3),
      pl_clk2 => ps_out.FCLK(2),
      pl_clk1 => ps_out.FCLK(1),
      pl_clk0 => ps_out.FCLK(0),

--------------------------
-- ACE interface allotment
--------------------------
      sacefpd_awuser => (others => '0'), --[15:0]
      sacefpd_aruser => (others => '0'), --[15:0]

--Debug and Test signals
      test_adc_clk => (others => '0'), --[3:0]
      test_adc_in => (others => '0'), --[31:0]
      test_adc2_in => (others => '0'), --[31:0]
      test_db => open, --[15:0]
      test_adc_out => open, --[19:0]
      test_ams_osc => open, --[7:0]
      test_mon_data => open, --[15:0]
      test_dclk => '0',
      test_den => '0',
      test_dwe => '0',
      test_daddr => (others => '0'), --[7:0]
      test_di => (others => '0'), --[15:0]
      test_drdy => open,
      test_do => open, --[15:0]
      test_convst => '0',
      pstp_pl_clk => (others => '0'), --[3:0]
      pstp_pl_in => (others => '0'), --[31:0]
      pstp_pl_out => open, --[31:0]
      pstp_pl_ts => (others => '0'), --[31:0]
      fmio_test_gem_scanmux_1 => '0',
      fmio_test_gem_scanmux_2 => '0',
      test_char_mode_fpd_n => '0',
      test_char_mode_lpd_n => '0',
      fmio_test_io_char_scan_clock => '0',
      fmio_test_io_char_scanenable => '0',
      fmio_test_io_char_scan_in => '0',
      fmio_test_io_char_scan_out => open,
      fmio_test_io_char_scan_reset_n => '0',
      fmio_char_afifslpd_test_select_n => '0',
      fmio_char_afifslpd_test_input => '0',
      fmio_char_afifslpd_test_output => open,
      fmio_char_afifsfpd_test_select_n => '0',
      fmio_char_afifsfpd_test_input => '0',
      fmio_char_afifsfpd_test_output => open,
      io_char_audio_in_test_data => '0',
      io_char_audio_mux_sel_n => '0',
      io_char_video_in_test_data => '0',
      io_char_video_mux_sel_n => '0',
      io_char_video_out_test_data => open,
      io_char_audio_out_test_data => open,
      fmio_test_qspi_scanmux_1_n => '0',
      fmio_test_sdio_scanmux_1 => '0',
      fmio_test_sdio_scanmux_2 => '0',
      fmio_sd0_dll_test_in_n => (others => '0'), --[3:0]
      fmio_sd0_dll_test_out => open, --[7:0]
      fmio_sd1_dll_test_in_n => (others => '0'), --[3:0]
      fmio_sd1_dll_test_out => open, --[7:0]
      test_pl_scan_chopper_si => '0',
      test_pl_scan_chopper_so => open,
      test_pl_scan_chopper_trig => '0',
      test_pl_scan_clk0 => '0',
      test_pl_scan_clk1 => '0',
      test_pl_scan_edt_clk => '0',
      test_pl_scan_edt_in_apu => '0',
      test_pl_scan_edt_in_cpu => '0',
      test_pl_scan_edt_in_ddr => (others => '0'), --[3:0]
      test_pl_scan_edt_in_fp => (others => '0'), --[9:0]
      test_pl_scan_edt_in_gpu => (others => '0'), --[3:0]
      test_pl_scan_edt_in_lp => (others => '0'), --[8:0]
      test_pl_scan_edt_in_usb3 => (others => '0'), --[1:0]
      test_pl_scan_edt_out_apu => open,
      test_pl_scan_edt_out_cpu0 => open,
      test_pl_scan_edt_out_cpu1 => open,
      test_pl_scan_edt_out_cpu2 => open,
      test_pl_scan_edt_out_cpu3 => open,
      test_pl_scan_edt_out_ddr => open, --[3:0]
      test_pl_scan_edt_out_fp => open, --[9:0]
      test_pl_scan_edt_out_gpu => open, --[3:0]
      test_pl_scan_edt_out_lp => open, --[8:0]
      test_pl_scan_edt_out_usb3 => open, --[1:0]
      test_pl_scan_edt_update => '0',
      test_pl_scan_reset_n => '0',
      test_pl_scanenable => '0',
      test_pl_scan_pll_reset => '0',
      test_pl_scan_spare_in0 => '0',
      test_pl_scan_spare_in1 => '0',
      test_pl_scan_spare_out0 => open,
      test_pl_scan_spare_out1 => open,
      test_pl_scan_wrap_clk => '0',
      test_pl_scan_wrap_ishift => '0',
      test_pl_scan_wrap_oshift => '0',
      test_pl_scan_slcr_config_clk => '0',
      test_pl_scan_slcr_config_rstn => '0',
      test_pl_scan_slcr_config_si => '0',
      test_pl_scan_spare_in2 => '0',
      test_pl_scanenable_slcr_en => '0',
      test_pl_pll_lock_out => open, --[4:0]
      test_pl_scan_slcr_config_so => open,
      tst_rtc_calibreg_in => (others => '0'), --[20:0]
      tst_rtc_calibreg_out => open, --[20:0]
      tst_rtc_calibreg_we => '0',
      tst_rtc_clk => '0',
      tst_rtc_osc_clk_out => open,
      tst_rtc_sec_counter_out => open, --[31:0]
      tst_rtc_seconds_raw_int => open,
      tst_rtc_testclock_select_n => '0',
      tst_rtc_tick_counter_out => open, --[15:0]
      tst_rtc_timesetreg_in => (others => '0'), --[31:0]
      tst_rtc_timesetreg_out => open, --[31:0]
      tst_rtc_disable_bat_op => '0',
      tst_rtc_osc_cntrl_in => (others => '0'), --[3:0]
      tst_rtc_osc_cntrl_out => open, --[3:0]
      tst_rtc_osc_cntrl_we => '0',
      tst_rtc_sec_reload => '0',
      tst_rtc_timesetreg_we => '0',
      tst_rtc_testmode_n => '0',
      test_usb0_funcmux_0_n => '0',
      test_usb1_funcmux_0_n => '0',
      test_usb0_scanmux_0_n => '0',
      test_usb1_scanmux_0_n => '0',
      lpd_pll_test_out => open, --[31:0]
      pl_lpd_pll_test_ck_sel_n => (others => '0'), --[2:0]
      pl_lpd_pll_test_fract_clk_sel_n => '0',
      pl_lpd_pll_test_fract_en_n => '0',
      pl_lpd_pll_test_mux_sel => '0',
      pl_lpd_pll_test_sel => (others => '0'), --[3:0]
      fpd_pll_test_out => open, --[31:0]
      pl_fpd_pll_test_ck_sel_n => (others => '0'), --[2:0]
      pl_fpd_pll_test_fract_clk_sel_n => '0',
      pl_fpd_pll_test_fract_en_n => '0',
      pl_fpd_pll_test_mux_sel => (others => '0'), --[1:0]
      pl_fpd_pll_test_sel => (others => '0'), --[3:0]
      fmio_char_gem_selection => (others => '0'), --[1:0]
      fmio_char_gem_test_select_n => '0',
      fmio_char_gem_test_input => '0',
      fmio_char_gem_test_output => open,
      test_ddr2pl_dcd_skewout => open,
      test_pl2ddr_dcd_sample_pulse => '0',
      test_bscan_en_n => '0',
      test_bscan_tdi => '0',
      test_bscan_updatedr => '0',
      test_bscan_shiftdr => '0',
      test_bscan_reset_tap_b => '0',
      test_bscan_misr_jtag_load => '0',
      test_bscan_intest => '0',
      test_bscan_extest => '0',
      test_bscan_clockdr => '0',
      test_bscan_ac_mode => '0',
      test_bscan_ac_test => '0',
      test_bscan_init_memory => '0',
      test_bscan_mode_c => '0',
      test_bscan_tdo => open,
      i_dbg_l0_txclk => '0',
      i_dbg_l0_rxclk => '0',
      i_dbg_l1_txclk => '0',
      i_dbg_l1_rxclk => '0',
      i_dbg_l2_txclk => '0',
      i_dbg_l2_rxclk => '0',
      i_dbg_l3_txclk => '0',
      i_dbg_l3_rxclk => '0',
      i_afe_rx_symbol_clk_by_2_pl => '0',
      pl_fpd_spare_0_in => '0',
      pl_fpd_spare_1_in => '0',
      pl_fpd_spare_2_in => '0',
      pl_fpd_spare_3_in => '0',
      pl_fpd_spare_4_in => '0',
      fpd_pl_spare_0_out => open,
      fpd_pl_spare_1_out => open,
      fpd_pl_spare_2_out => open,
      fpd_pl_spare_3_out => open,
      fpd_pl_spare_4_out => open,
      pl_lpd_spare_0_in => '0',
      pl_lpd_spare_1_in => '0',
      pl_lpd_spare_2_in => '0',
      pl_lpd_spare_3_in => '0',
      pl_lpd_spare_4_in => '0',
      lpd_pl_spare_0_out => open,
      lpd_pl_spare_1_out => open,
      lpd_pl_spare_2_out => open,
      lpd_pl_spare_3_out => open,
      lpd_pl_spare_4_out => open,
      o_dbg_l0_phystatus => open,
      o_dbg_l0_rxdata => open, --[19:0]
      o_dbg_l0_rxdatak => open, --[1:0]
      o_dbg_l0_rxvalid => open,
      o_dbg_l0_rxstatus => open, --[2:0]
      o_dbg_l0_rxelecidle => open,
      o_dbg_l0_rstb => open,
      o_dbg_l0_txdata => open, --[19:0]
      o_dbg_l0_txdatak => open, --[1:0]
      o_dbg_l0_rate => open, --[1:0]
      o_dbg_l0_powerdown => open, --[1:0]
      o_dbg_l0_txelecidle => open,
      o_dbg_l0_txdetrx_lpback => open,
      o_dbg_l0_rxpolarity => open,
      o_dbg_l0_tx_sgmii_ewrap => open,
      o_dbg_l0_rx_sgmii_en_cdet => open,
      o_dbg_l0_sata_corerxdata => open, --[19:0]
      o_dbg_l0_sata_corerxdatavalid => open, --[1:0]
      o_dbg_l0_sata_coreready => open,
      o_dbg_l0_sata_coreclockready => open,
      o_dbg_l0_sata_corerxsignaldet => open,
      o_dbg_l0_sata_phyctrltxdata => open, --[19:0]
      o_dbg_l0_sata_phyctrltxidle => open,
      o_dbg_l0_sata_phyctrltxrate => open, --[1:0]
      o_dbg_l0_sata_phyctrlrxrate => open, --[1:0]
      o_dbg_l0_sata_phyctrltxrst => open,
      o_dbg_l0_sata_phyctrlrxrst => open,
      o_dbg_l0_sata_phyctrlreset => open,
      o_dbg_l0_sata_phyctrlpartial => open,
      o_dbg_l0_sata_phyctrlslumber => open,
      o_dbg_l1_phystatus => open,
      o_dbg_l1_rxdata => open, --[19:0]
      o_dbg_l1_rxdatak => open, --[1:0]
      o_dbg_l1_rxvalid => open,
      o_dbg_l1_rxstatus => open, --[2:0]
      o_dbg_l1_rxelecidle => open,
      o_dbg_l1_rstb => open,
      o_dbg_l1_txdata => open, --[19:0]
      o_dbg_l1_txdatak => open, --[1:0]
      o_dbg_l1_rate => open, --[1:0]
      o_dbg_l1_powerdown => open, --[1:0]
      o_dbg_l1_txelecidle => open,
      o_dbg_l1_txdetrx_lpback => open,
      o_dbg_l1_rxpolarity => open,
      o_dbg_l1_tx_sgmii_ewrap => open,
      o_dbg_l1_rx_sgmii_en_cdet => open,
      o_dbg_l1_sata_corerxdata => open, --[19:0]
      o_dbg_l1_sata_corerxdatavalid => open, --[1:0]
      o_dbg_l1_sata_coreready => open,
      o_dbg_l1_sata_coreclockready => open,
      o_dbg_l1_sata_corerxsignaldet => open,
      o_dbg_l1_sata_phyctrltxdata => open, --[19:0]
      o_dbg_l1_sata_phyctrltxidle => open,
      o_dbg_l1_sata_phyctrltxrate => open, --[1:0]
      o_dbg_l1_sata_phyctrlrxrate => open, --[1:0]
      o_dbg_l1_sata_phyctrltxrst => open,
      o_dbg_l1_sata_phyctrlrxrst => open,
      o_dbg_l1_sata_phyctrlreset => open,
      o_dbg_l1_sata_phyctrlpartial => open,
      o_dbg_l1_sata_phyctrlslumber => open,
      o_dbg_l2_phystatus => open,
      o_dbg_l2_rxdata => open, --[19:0]
      o_dbg_l2_rxdatak => open, --[1:0]
      o_dbg_l2_rxvalid => open,
      o_dbg_l2_rxstatus => open, --[2:0]
      o_dbg_l2_rxelecidle => open,
      o_dbg_l2_rstb => open,
      o_dbg_l2_txdata => open, --[19:0]
      o_dbg_l2_txdatak => open, --[1:0]
      o_dbg_l2_rate => open, --[1:0]
      o_dbg_l2_powerdown => open, --[1:0]
      o_dbg_l2_txelecidle => open,
      o_dbg_l2_txdetrx_lpback => open,
      o_dbg_l2_rxpolarity => open,
      o_dbg_l2_tx_sgmii_ewrap => open,
      o_dbg_l2_rx_sgmii_en_cdet => open,
      o_dbg_l2_sata_corerxdata => open, --[19:0]
      o_dbg_l2_sata_corerxdatavalid => open, --[1:0]
      o_dbg_l2_sata_coreready => open,
      o_dbg_l2_sata_coreclockready => open,
      o_dbg_l2_sata_corerxsignaldet => open,
      o_dbg_l2_sata_phyctrltxdata => open, --[19:0]
      o_dbg_l2_sata_phyctrltxidle => open,
      o_dbg_l2_sata_phyctrltxrate => open, --[1:0]
      o_dbg_l2_sata_phyctrlrxrate => open, --[1:0]
      o_dbg_l2_sata_phyctrltxrst => open,
      o_dbg_l2_sata_phyctrlrxrst => open,
      o_dbg_l2_sata_phyctrlreset => open,
      o_dbg_l2_sata_phyctrlpartial => open,
      o_dbg_l2_sata_phyctrlslumber => open,
      o_dbg_l3_phystatus => open,
      o_dbg_l3_rxdata => open, --[19:0]
      o_dbg_l3_rxdatak => open, --[1:0]
      o_dbg_l3_rxvalid => open,
      o_dbg_l3_rxstatus => open, --[2:0]
      o_dbg_l3_rxelecidle => open,
      o_dbg_l3_rstb => open,
      o_dbg_l3_txdata => open, --[19:0]
      o_dbg_l3_txdatak => open, --[1:0]
      o_dbg_l3_rate => open, --[1:0]
      o_dbg_l3_powerdown => open, --[1:0]
      o_dbg_l3_txelecidle => open,
      o_dbg_l3_txdetrx_lpback => open,
      o_dbg_l3_rxpolarity => open,
      o_dbg_l3_tx_sgmii_ewrap => open,
      o_dbg_l3_rx_sgmii_en_cdet => open,
      o_dbg_l3_sata_corerxdata => open, --[19:0]
      o_dbg_l3_sata_corerxdatavalid => open, --[1:0]
      o_dbg_l3_sata_coreready => open,
      o_dbg_l3_sata_coreclockready => open,
      o_dbg_l3_sata_corerxsignaldet => open,
      o_dbg_l3_sata_phyctrltxdata => open, --[19:0]
      o_dbg_l3_sata_phyctrltxidle => open,
      o_dbg_l3_sata_phyctrltxrate => open, --[1:0]
      o_dbg_l3_sata_phyctrlrxrate => open, --[1:0]
      o_dbg_l3_sata_phyctrltxrst => open,
      o_dbg_l3_sata_phyctrlrxrst => open,
      o_dbg_l3_sata_phyctrlreset => open,
      o_dbg_l3_sata_phyctrlpartial => open,
      o_dbg_l3_sata_phyctrlslumber => open,
      dbg_path_fifo_bypass => open,
      i_afe_pll_pd_hs_clock_r => '0',
      i_afe_mode => '0',
      i_bgcal_afe_mode => '0',
      o_afe_cmn_calib_comp_out => open,
      i_afe_cmn_bg_enable_low_leakage => '0',
      i_afe_cmn_bg_iso_ctrl_bar => '0',
      i_afe_cmn_bg_pd => '0',
      i_afe_cmn_bg_pd_bg_ok => '0',
      i_afe_cmn_bg_pd_ptat => '0',
      i_afe_cmn_calib_en_iconst => '0',
      i_afe_cmn_calib_enable_low_leakage => '0',
      i_afe_cmn_calib_iso_ctrl_bar => '0',
      o_afe_pll_dco_count => open, --[12:0]
      o_afe_pll_clk_sym_hs => open,
      o_afe_pll_fbclk_frac => open,
      o_afe_rx_pipe_lfpsbcn_rxelecidle => open,
      o_afe_rx_pipe_sigdet => open,
      o_afe_rx_symbol => open, --[19:0]
      o_afe_rx_symbol_clk_by_2 => open,
      o_afe_rx_uphy_save_calcode => open,
      o_afe_rx_uphy_startloop_buf => open,
      o_afe_rx_uphy_rx_calib_done => open,
      i_afe_rx_rxpma_rstb => '0',
      i_afe_rx_uphy_restore_calcode_data => (others => '0'), --[7:0]
      i_afe_rx_pipe_rxeqtraining => '0',
      i_afe_rx_iso_hsrx_ctrl_bar => '0',
      i_afe_rx_iso_lfps_ctrl_bar => '0',
      i_afe_rx_iso_sigdet_ctrl_bar => '0',
      i_afe_rx_hsrx_clock_stop_req => '0',
      o_afe_rx_uphy_save_calcode_data => open, --[7:0]
      o_afe_rx_hsrx_clock_stop_ack => open,
      o_afe_pg_avddcr => open,
      o_afe_pg_avddio => open,
      o_afe_pg_dvddcr => open,
      o_afe_pg_static_avddcr => open,
      o_afe_pg_static_avddio => open,
      i_pll_afe_mode => '0',
      i_afe_pll_coarse_code => (others => '0'), --[10:0]
      i_afe_pll_en_clock_hs_div2 => '0',
      i_afe_pll_fbdiv => (others => '0'), --[15:0]
      i_afe_pll_load_fbdiv => '0',
      i_afe_pll_pd => '0',
      i_afe_pll_pd_pfd => '0',
      i_afe_pll_rst_fdbk_div => '0',
      i_afe_pll_startloop => '0',
      i_afe_pll_v2i_code => (others => '0'), --[5:0]
      i_afe_pll_v2i_prog => (others => '0'), --[4:0]
      i_afe_pll_vco_cnt_window => '0',
      i_afe_rx_mphy_gate_symbol_clk => '0',
      i_afe_rx_mphy_mux_hsb_ls => '0',
      i_afe_rx_pipe_rx_term_enable => '0',
      i_afe_rx_uphy_biasgen_iconst_core_mirror_enable => '0',
      i_afe_rx_uphy_biasgen_iconst_io_mirror_enable => '0',
      i_afe_rx_uphy_biasgen_irconst_core_mirror_enable => '0',
      i_afe_rx_uphy_enable_cdr => '0',
      i_afe_rx_uphy_enable_low_leakage => '0',
      i_afe_rx_rxpma_refclk_dig => '0',
      i_afe_rx_uphy_hsrx_rstb => '0',
      i_afe_rx_uphy_pdn_hs_des => '0',
      i_afe_rx_uphy_pd_samp_c2c => '0',
      i_afe_rx_uphy_pd_samp_c2c_eclk => '0',
      i_afe_rx_uphy_pso_clk_lane => '0',
      i_afe_rx_uphy_pso_eq => '0',
      i_afe_rx_uphy_pso_hsrxdig => '0',
      i_afe_rx_uphy_pso_iqpi => '0',
      i_afe_rx_uphy_pso_lfpsbcn => '0',
      i_afe_rx_uphy_pso_samp_flops => '0',
      i_afe_rx_uphy_pso_sigdet => '0',
      i_afe_rx_uphy_restore_calcode => '0',
      i_afe_rx_uphy_run_calib => '0',
      i_afe_rx_uphy_rx_lane_polarity_swap => '0',
      i_afe_rx_uphy_startloop_pll => '0',
      i_afe_rx_uphy_hsclk_division_factor => (others => '0'), --[1:0]
      i_afe_rx_uphy_rx_pma_opmode => (others => '0'), --[7:0]
      i_afe_tx_enable_hsclk_division => (others => '0'), --[1:0]
      i_afe_tx_enable_ldo => '0',
      i_afe_tx_enable_ref => '0',
      i_afe_tx_enable_supply_hsclk => '0',
      i_afe_tx_enable_supply_pipe => '0',
      i_afe_tx_enable_supply_serializer => '0',
      i_afe_tx_enable_supply_uphy => '0',
      i_afe_tx_hs_ser_rstb => '0',
      i_afe_tx_hs_symbol => (others => '0'), --[19:0]
      i_afe_tx_mphy_tx_ls_data => '0',
      i_afe_tx_pipe_tx_enable_idle_mode => (others => '0'), --[1:0]
      i_afe_tx_pipe_tx_enable_lfps => (others => '0'), --[1:0]
      i_afe_tx_pipe_tx_enable_rxdet => '0',
      i_afe_TX_uphy_txpma_opmode => (others => '0'), --[7:0]
      i_afe_TX_pmadig_digital_reset_n => '0',
      i_afe_TX_serializer_rst_rel => '0',
      i_afe_TX_pll_symb_clk_2 => '0',
      i_afe_TX_ana_if_rate => (others => '0'), --[1:0]
      i_afe_TX_en_dig_sublp_mode => '0',
      i_afe_TX_LPBK_SEL => (others => '0'), --[2:0]
      i_afe_TX_iso_ctrl_bar => '0',
      i_afe_TX_ser_iso_ctrl_bar => '0',
      i_afe_TX_lfps_clk => '0',
      i_afe_TX_serializer_rstb => '0',
      o_afe_TX_dig_reset_rel_ack => open,
      o_afe_TX_pipe_TX_dn_rxdet => open,
      o_afe_TX_pipe_TX_dp_rxdet => open,
      i_afe_tx_pipe_tx_fast_est_common_mode => '0',
      o_dbg_l0_txclk => open,
      o_dbg_l0_rxclk => open,
      o_dbg_l1_txclk => open,
      o_dbg_l1_rxclk => open,
      o_dbg_l2_txclk => open,
      o_dbg_l2_rxclk => open,
      o_dbg_l3_txclk => open,
      o_dbg_l3_rxclk => open
      );
end rtl;
