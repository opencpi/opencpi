-- THIS FILE WAS ORIGINALLY GENERATED ON Thu Aug 30 20:34:00 2012 EDT
-- BASED ON THE FILE: sym_fir_real.xml
-- YOU ARE EXPECTED TO EDIT IT
-- This file contains the architecture skeleton for worker: sym_fir_real

library IEEE;
  use IEEE.std_logic_1164.all;

architecture rtl of sym_fir_real is
begin -- rtl



end rtl;
