../../../comparator_real.rcc/target-macos-10_9-x86_64/generics.vhd