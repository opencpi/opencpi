../../../file_write_msg.rcc/target-linux-c6-x86_64/generics.vhd