// THIS FILE WAS ORIGINALLY GENERATED ON Thu Sep 20 16:26:19 2012 EDT
// BASED ON THE FILE: fft1d.xml
// YOU ARE EXPECTED TO EDIT IT
// This file contains the implementation skeleton for worker: fft1d

`include "fft1d-impl.vh"



endmodule //fft1d
