// Hand Edited from generated verilog to:
// 1. Move config ROM outside this module since can change after this is synthesized...
// 2. Move time server outside this module since it might be platform-specific and is not "CP".
// 3. Move DNA outside this module since it is platform-specific.
// 4. UUID and ROM are moved elsewhere entirely
// 5. PCIdevice is moved elsewhere
//
// Notes about fixing the fact that the BSV master side is not doing the OK and Error responses,
// but only the timeout and reset responses.
// Master: Checks for failure, but always copies the response data.
// Need to identify the entry to the response FIFO
// MUX_wci_respF{_N}$enq_1__VAL_1 looks like the load value
// Others are _VAL_2,3,4,5,6,7
// Val_1: if resp is null, timeout, else response: used on SEL_1
// Val_2: wci_wStatus: used on      WILL_FIRE_RL_cpDispatch_F_F_F_F_T_F_F_T:
// Val_3: x_data__h104757 : used on WILL_FIRE_RL_cpDispatch_F_F_F_F_T_F_F_F_T:
//          reset and control register
// Val_4: x_data__h104763 : used on WILL_FIRE_RL_cpDispatch_F_F_F_F_T_F_F_F_F_T:
//          last config addr
// Val_5: pagewindow : used on      WILL_FIRE_RL_cpDispatch_F_F_F_F_T_F_F_F_F_F_T:
// 34'h100000000: used on           MUX_wci_respF$enq_1__SEL_6
//       Ack of control write
// 34'h1C0DE4204; used on           MUX_wci_respF$enq_1__SEL_7
//       RESET error
// 34'h3C0DE4202; used on           WILL_FIRE_RL_cpDispatch_F_F_T_T_F_T:
//       Worker ERROR on control op write
// Generated by Bluespec Compiler, version 2012.09.beta1 (build 29570, 2012-09.11)
//
// On Wed Oct 24 10:26:52 EDT 2012
//
//
// Ports:
// Name                         I/O  size props
// RDY_server_request_put         O     1 reg
// server_response_get            O    40 reg
// RDY_server_response_get        O     1 reg
// wci_Vm_0_MCmd                  O     3
// wci_Vm_0_MAddrSpace            O     1
// wci_Vm_0_MByteEn               O     4
// wci_Vm_0_MAddr                 O    32
// wci_Vm_0_MData                 O    32 reg
// wci_Vm_0_MFlag                 O     2 reg
// wci_Vm_1_MCmd                  O     3
// wci_Vm_1_MAddrSpace            O     1
// wci_Vm_1_MByteEn               O     4
// wci_Vm_1_MAddr                 O    32
// wci_Vm_1_MData                 O    32 reg
// wci_Vm_1_MFlag                 O     2 reg
// wci_Vm_2_MCmd                  O     3
// wci_Vm_2_MAddrSpace            O     1
// wci_Vm_2_MByteEn               O     4
// wci_Vm_2_MAddr                 O    32
// wci_Vm_2_MData                 O    32 reg
// wci_Vm_2_MFlag                 O     2 reg
// wci_Vm_3_MCmd                  O     3
// wci_Vm_3_MAddrSpace            O     1
// wci_Vm_3_MByteEn               O     4
// wci_Vm_3_MAddr                 O    32
// wci_Vm_3_MData                 O    32 reg
// wci_Vm_3_MFlag                 O     2 reg
// wci_Vm_4_MCmd                  O     3
// wci_Vm_4_MAddrSpace            O     1
// wci_Vm_4_MByteEn               O     4
// wci_Vm_4_MAddr                 O    32
// wci_Vm_4_MData                 O    32 reg
// wci_Vm_4_MFlag                 O     2 reg
// wci_Vm_5_MCmd                  O     3
// wci_Vm_5_MAddrSpace            O     1
// wci_Vm_5_MByteEn               O     4
// wci_Vm_5_MAddr                 O    32
// wci_Vm_5_MData                 O    32 reg
// wci_Vm_5_MFlag                 O     2 reg
// wci_Vm_6_MCmd                  O     3
// wci_Vm_6_MAddrSpace            O     1
// wci_Vm_6_MByteEn               O     4
// wci_Vm_6_MAddr                 O    32
// wci_Vm_6_MData                 O    32 reg
// wci_Vm_6_MFlag                 O     2 reg
// wci_Vm_7_MCmd                  O     3
// wci_Vm_7_MAddrSpace            O     1
// wci_Vm_7_MByteEn               O     4
// wci_Vm_7_MAddr                 O    32
// wci_Vm_7_MData                 O    32 reg
// wci_Vm_7_MFlag                 O     2 reg
// wci_Vm_8_MCmd                  O     3
// wci_Vm_8_MAddrSpace            O     1
// wci_Vm_8_MByteEn               O     4
// wci_Vm_8_MAddr                 O    32
// wci_Vm_8_MData                 O    32 reg
// wci_Vm_8_MFlag                 O     2 reg
// wci_Vm_9_MCmd                  O     3
// wci_Vm_9_MAddrSpace            O     1
// wci_Vm_9_MByteEn               O     4
// wci_Vm_9_MAddr                 O    32
// wci_Vm_9_MData                 O    32 reg
// wci_Vm_9_MFlag                 O     2 reg
// wci_Vm_10_MCmd                 O     3
// wci_Vm_10_MAddrSpace           O     1
// wci_Vm_10_MByteEn              O     4
// wci_Vm_10_MAddr                O    32
// wci_Vm_10_MData                O    32 reg
// wci_Vm_10_MFlag                O     2 reg
// wci_Vm_11_MCmd                 O     3
// wci_Vm_11_MAddrSpace           O     1
// wci_Vm_11_MByteEn              O     4
// wci_Vm_11_MAddr                O    32
// wci_Vm_11_MData                O    32 reg
// wci_Vm_11_MFlag                O     2 reg
// wci_Vm_12_MCmd                 O     3
// wci_Vm_12_MAddrSpace           O     1
// wci_Vm_12_MByteEn              O     4
// wci_Vm_12_MAddr                O    32
// wci_Vm_12_MData                O    32 reg
// wci_Vm_12_MFlag                O     2 reg
// wci_Vm_13_MCmd                 O     3
// wci_Vm_13_MAddrSpace           O     1
// wci_Vm_13_MByteEn              O     4
// wci_Vm_13_MAddr                O    32
// wci_Vm_13_MData                O    32 reg
// wci_Vm_13_MFlag                O     2 reg
// wci_Vm_14_MCmd                 O     3
// wci_Vm_14_MAddrSpace           O     1
// wci_Vm_14_MByteEn              O     4
// wci_Vm_14_MAddr                O    32
// wci_Vm_14_MData                O    32 reg
// wci_Vm_14_MFlag                O     2 reg
// cpNow                          O    64 reg
// RDY_cpNow                      O     1 const
// gps_ppsSyncOut                 O     1
// led                            O     2 reg
// RST_N_wci_Vm_0                 O     1 reset
// RST_N_wci_Vm_1                 O     1 reset
// RST_N_wci_Vm_2                 O     1 reset
// RST_N_wci_Vm_3                 O     1 reset
// RST_N_wci_Vm_4                 O     1 reset
// RST_N_wci_Vm_5                 O     1 reset
// RST_N_wci_Vm_6                 O     1 reset
// RST_N_wci_Vm_7                 O     1 reset
// RST_N_wci_Vm_8                 O     1 reset
// RST_N_wci_Vm_9                 O     1 reset
// RST_N_wci_Vm_10                O     1 reset
// RST_N_wci_Vm_11                O     1 reset
// RST_N_wci_Vm_12                O     1 reset
// RST_N_wci_Vm_13                O     1 reset
// RST_N_wci_Vm_14                O     1 reset
// pciDevice                      I    16
// CLK_time_clk                   I     1 clock
// RST_N_time_rst                 I     1 reset
// CLK                            I     1 clock
// RST_N                          I     1 reset
// server_request_put             I    59 reg
// wci_Vm_0_SResp                 I     2
// wci_Vm_0_SData                 I    32
// wci_Vm_0_SFlag                 I     2 reg
// wci_Vm_1_SResp                 I     2
// wci_Vm_1_SData                 I    32
// wci_Vm_1_SFlag                 I     2 reg
// wci_Vm_2_SResp                 I     2
// wci_Vm_2_SData                 I    32
// wci_Vm_2_SFlag                 I     2 reg
// wci_Vm_3_SResp                 I     2
// wci_Vm_3_SData                 I    32
// wci_Vm_3_SFlag                 I     2 reg
// wci_Vm_4_SResp                 I     2
// wci_Vm_4_SData                 I    32
// wci_Vm_4_SFlag                 I     2 reg
// wci_Vm_5_SResp                 I     2
// wci_Vm_5_SData                 I    32
// wci_Vm_5_SFlag                 I     2 reg
// wci_Vm_6_SResp                 I     2
// wci_Vm_6_SData                 I    32
// wci_Vm_6_SFlag                 I     2 reg
// wci_Vm_7_SResp                 I     2
// wci_Vm_7_SData                 I    32
// wci_Vm_7_SFlag                 I     2 reg
// wci_Vm_8_SResp                 I     2
// wci_Vm_8_SData                 I    32
// wci_Vm_8_SFlag                 I     2 reg
// wci_Vm_9_SResp                 I     2
// wci_Vm_9_SData                 I    32
// wci_Vm_9_SFlag                 I     2 reg
// wci_Vm_10_SResp                I     2
// wci_Vm_10_SData                I    32
// wci_Vm_10_SFlag                I     2 reg
// wci_Vm_11_SResp                I     2
// wci_Vm_11_SData                I    32
// wci_Vm_11_SFlag                I     2 reg
// wci_Vm_12_SResp                I     2
// wci_Vm_12_SData                I    32
// wci_Vm_12_SFlag                I     2 reg
// wci_Vm_13_SResp                I     2
// wci_Vm_13_SData                I    32
// wci_Vm_13_SFlag                I     2 reg
// wci_Vm_14_SResp                I     2
// wci_Vm_14_SData                I    32
// wci_Vm_14_SFlag                I     2 reg
// gps_ppsSyncIn_x                I     1 reg
// switch_x                       I     3 reg
// uuid_arg                       I   512
// EN_server_request_put          I     1
// wci_Vm_0_SThreadBusy           I     1 reg
// wci_Vm_1_SThreadBusy           I     1 reg
// wci_Vm_2_SThreadBusy           I     1 reg
// wci_Vm_3_SThreadBusy           I     1 reg
// wci_Vm_4_SThreadBusy           I     1 reg
// wci_Vm_5_SThreadBusy           I     1 reg
// wci_Vm_6_SThreadBusy           I     1 reg
// wci_Vm_7_SThreadBusy           I     1 reg
// wci_Vm_8_SThreadBusy           I     1 reg
// wci_Vm_9_SThreadBusy           I     1 reg
// wci_Vm_10_SThreadBusy          I     1 reg
// wci_Vm_11_SThreadBusy          I     1 reg
// wci_Vm_12_SThreadBusy          I     1 reg
// wci_Vm_13_SThreadBusy          I     1 reg
// wci_Vm_14_SThreadBusy          I     1 reg
// EN_server_response_get         I     1
//
// No combinational paths from inputs to outputs
//
//

`ifdef BSV_ASSIGNMENT_DELAY
`else
  `define BSV_ASSIGNMENT_DELAY
`endif

`ifdef BSV_POSITIVE_RESET
  `define BSV_RESET_VALUE 1'b1
  `define BSV_RESET_EDGE posedge
`else
  `define BSV_RESET_VALUE 1'b0
  `define BSV_RESET_EDGE negedge
`endif

`ifdef not
module mkOCCP(pciDevice,
	      CLK_time_clk,
	      RST_N_time_rst,
`else
module mkOCCP(
`endif
	      CLK,
	      RST_N,

	      server_request_put,
	      EN_server_request_put,
	      RDY_server_request_put,

	      EN_server_response_get,
	      server_response_get,
	      RDY_server_response_get,

	      wci_Vm_0_MCmd,

	      wci_Vm_0_MAddrSpace,

	      wci_Vm_0_MByteEn,

	      wci_Vm_0_MAddr,

	      wci_Vm_0_MData,

	      wci_Vm_0_SResp,

	      wci_Vm_0_SData,

	      wci_Vm_0_SThreadBusy,

	      wci_Vm_0_SFlag,

	      wci_Vm_0_MFlag,

	      wci_Vm_1_MCmd,

	      wci_Vm_1_MAddrSpace,

	      wci_Vm_1_MByteEn,

	      wci_Vm_1_MAddr,

	      wci_Vm_1_MData,

	      wci_Vm_1_SResp,

	      wci_Vm_1_SData,

	      wci_Vm_1_SThreadBusy,

	      wci_Vm_1_SFlag,

	      wci_Vm_1_MFlag,

	      wci_Vm_2_MCmd,

	      wci_Vm_2_MAddrSpace,

	      wci_Vm_2_MByteEn,

	      wci_Vm_2_MAddr,

	      wci_Vm_2_MData,

	      wci_Vm_2_SResp,

	      wci_Vm_2_SData,

	      wci_Vm_2_SThreadBusy,

	      wci_Vm_2_SFlag,

	      wci_Vm_2_MFlag,

	      wci_Vm_3_MCmd,

	      wci_Vm_3_MAddrSpace,

	      wci_Vm_3_MByteEn,

	      wci_Vm_3_MAddr,

	      wci_Vm_3_MData,

	      wci_Vm_3_SResp,

	      wci_Vm_3_SData,

	      wci_Vm_3_SThreadBusy,

	      wci_Vm_3_SFlag,

	      wci_Vm_3_MFlag,

	      wci_Vm_4_MCmd,

	      wci_Vm_4_MAddrSpace,

	      wci_Vm_4_MByteEn,

	      wci_Vm_4_MAddr,

	      wci_Vm_4_MData,

	      wci_Vm_4_SResp,

	      wci_Vm_4_SData,

	      wci_Vm_4_SThreadBusy,

	      wci_Vm_4_SFlag,

	      wci_Vm_4_MFlag,

	      wci_Vm_5_MCmd,

	      wci_Vm_5_MAddrSpace,

	      wci_Vm_5_MByteEn,

	      wci_Vm_5_MAddr,

	      wci_Vm_5_MData,

	      wci_Vm_5_SResp,

	      wci_Vm_5_SData,

	      wci_Vm_5_SThreadBusy,

	      wci_Vm_5_SFlag,

	      wci_Vm_5_MFlag,

	      wci_Vm_6_MCmd,

	      wci_Vm_6_MAddrSpace,

	      wci_Vm_6_MByteEn,

	      wci_Vm_6_MAddr,

	      wci_Vm_6_MData,

	      wci_Vm_6_SResp,

	      wci_Vm_6_SData,

	      wci_Vm_6_SThreadBusy,

	      wci_Vm_6_SFlag,

	      wci_Vm_6_MFlag,

	      wci_Vm_7_MCmd,

	      wci_Vm_7_MAddrSpace,

	      wci_Vm_7_MByteEn,

	      wci_Vm_7_MAddr,

	      wci_Vm_7_MData,

	      wci_Vm_7_SResp,

	      wci_Vm_7_SData,

	      wci_Vm_7_SThreadBusy,

	      wci_Vm_7_SFlag,

	      wci_Vm_7_MFlag,

	      wci_Vm_8_MCmd,

	      wci_Vm_8_MAddrSpace,

	      wci_Vm_8_MByteEn,

	      wci_Vm_8_MAddr,

	      wci_Vm_8_MData,

	      wci_Vm_8_SResp,

	      wci_Vm_8_SData,

	      wci_Vm_8_SThreadBusy,

	      wci_Vm_8_SFlag,

	      wci_Vm_8_MFlag,

	      wci_Vm_9_MCmd,

	      wci_Vm_9_MAddrSpace,

	      wci_Vm_9_MByteEn,

	      wci_Vm_9_MAddr,

	      wci_Vm_9_MData,

	      wci_Vm_9_SResp,

	      wci_Vm_9_SData,

	      wci_Vm_9_SThreadBusy,

	      wci_Vm_9_SFlag,

	      wci_Vm_9_MFlag,

	      wci_Vm_10_MCmd,

	      wci_Vm_10_MAddrSpace,

	      wci_Vm_10_MByteEn,

	      wci_Vm_10_MAddr,

	      wci_Vm_10_MData,

	      wci_Vm_10_SResp,

	      wci_Vm_10_SData,

	      wci_Vm_10_SThreadBusy,

	      wci_Vm_10_SFlag,

	      wci_Vm_10_MFlag,

	      wci_Vm_11_MCmd,

	      wci_Vm_11_MAddrSpace,

	      wci_Vm_11_MByteEn,

	      wci_Vm_11_MAddr,

	      wci_Vm_11_MData,

	      wci_Vm_11_SResp,

	      wci_Vm_11_SData,

	      wci_Vm_11_SThreadBusy,

	      wci_Vm_11_SFlag,

	      wci_Vm_11_MFlag,

	      wci_Vm_12_MCmd,

	      wci_Vm_12_MAddrSpace,

	      wci_Vm_12_MByteEn,

	      wci_Vm_12_MAddr,

	      wci_Vm_12_MData,

	      wci_Vm_12_SResp,

	      wci_Vm_12_SData,

	      wci_Vm_12_SThreadBusy,

	      wci_Vm_12_SFlag,

	      wci_Vm_12_MFlag,

	      wci_Vm_13_MCmd,

	      wci_Vm_13_MAddrSpace,

	      wci_Vm_13_MByteEn,

	      wci_Vm_13_MAddr,

	      wci_Vm_13_MData,

	      wci_Vm_13_SResp,

	      wci_Vm_13_SData,

	      wci_Vm_13_SThreadBusy,

	      wci_Vm_13_SFlag,

	      wci_Vm_13_MFlag,

	      wci_Vm_14_MCmd,

	      wci_Vm_14_MAddrSpace,

	      wci_Vm_14_MByteEn,

	      wci_Vm_14_MAddr,

	      wci_Vm_14_MData,

	      wci_Vm_14_SResp,

	      wci_Vm_14_SData,

	      wci_Vm_14_SThreadBusy,

	      wci_Vm_14_SFlag,

	      wci_Vm_14_MFlag,

`ifdef not
	      cpNow,
	      RDY_cpNow,

	      gps_ppsSyncIn_x,

	      gps_ppsSyncOut,

	      led,

	      switch_x,

	      uuid_arg,
	      rom_en,
	      rom_addr,
	      rom_data,
`endif
	      
	      RST_N_wci_Vm_0,
	      RST_N_wci_Vm_1,
	      RST_N_wci_Vm_2,
	      RST_N_wci_Vm_3,
	      RST_N_wci_Vm_4,
	      RST_N_wci_Vm_5,
	      RST_N_wci_Vm_6,
	      RST_N_wci_Vm_7,
	      RST_N_wci_Vm_8,
	      RST_N_wci_Vm_9,
	      RST_N_wci_Vm_10,
	      RST_N_wci_Vm_11,
	      RST_N_wci_Vm_12,
	      RST_N_wci_Vm_13,
	      RST_N_wci_Vm_14);
`ifdef not
  input  [15 : 0] pciDevice;
  input  CLK_time_clk;
  input  RST_N_time_rst;
`endif
  input  CLK;
  input  RST_N;

  // action method server_request_put
  input  [58 : 0] server_request_put;
  input  EN_server_request_put;
  output RDY_server_request_put;

  // actionvalue method server_response_get
  input  EN_server_response_get;
  output [39 : 0] server_response_get;
  output RDY_server_response_get;

  // value method wci_Vm_0_mCmd
  output [2 : 0] wci_Vm_0_MCmd;

  // value method wci_Vm_0_mAddrSpace
  output wci_Vm_0_MAddrSpace;

  // value method wci_Vm_0_mByteEn
  output [3 : 0] wci_Vm_0_MByteEn;

  // value method wci_Vm_0_mAddr
  output [31 : 0] wci_Vm_0_MAddr;

  // value method wci_Vm_0_mData
  output [31 : 0] wci_Vm_0_MData;

  // action method wci_Vm_0_sResp
  input  [1 : 0] wci_Vm_0_SResp;

  // action method wci_Vm_0_sData
  input  [31 : 0] wci_Vm_0_SData;

  // action method wci_Vm_0_sThreadBusy
  input  wci_Vm_0_SThreadBusy;

  // action method wci_Vm_0_sFlag
  input  [2 : 0] wci_Vm_0_SFlag;

  // value method wci_Vm_0_mFlag
  output [1 : 0] wci_Vm_0_MFlag;

  // value method wci_Vm_1_mCmd
  output [2 : 0] wci_Vm_1_MCmd;

  // value method wci_Vm_1_mAddrSpace
  output wci_Vm_1_MAddrSpace;

  // value method wci_Vm_1_mByteEn
  output [3 : 0] wci_Vm_1_MByteEn;

  // value method wci_Vm_1_mAddr
  output [31 : 0] wci_Vm_1_MAddr;

  // value method wci_Vm_1_mData
  output [31 : 0] wci_Vm_1_MData;

  // action method wci_Vm_1_sResp
  input  [1 : 0] wci_Vm_1_SResp;

  // action method wci_Vm_1_sData
  input  [31 : 0] wci_Vm_1_SData;

  // action method wci_Vm_1_sThreadBusy
  input  wci_Vm_1_SThreadBusy;

  // action method wci_Vm_1_sFlag
  input  [2 : 0] wci_Vm_1_SFlag;

  // value method wci_Vm_1_mFlag
  output [1 : 0] wci_Vm_1_MFlag;

  // value method wci_Vm_2_mCmd
  output [2 : 0] wci_Vm_2_MCmd;

  // value method wci_Vm_2_mAddrSpace
  output wci_Vm_2_MAddrSpace;

  // value method wci_Vm_2_mByteEn
  output [3 : 0] wci_Vm_2_MByteEn;

  // value method wci_Vm_2_mAddr
  output [31 : 0] wci_Vm_2_MAddr;

  // value method wci_Vm_2_mData
  output [31 : 0] wci_Vm_2_MData;

  // action method wci_Vm_2_sResp
  input  [1 : 0] wci_Vm_2_SResp;

  // action method wci_Vm_2_sData
  input  [31 : 0] wci_Vm_2_SData;

  // action method wci_Vm_2_sThreadBusy
  input  wci_Vm_2_SThreadBusy;

  // action method wci_Vm_2_sFlag
  input  [2 : 0] wci_Vm_2_SFlag;

  // value method wci_Vm_2_mFlag
  output [1 : 0] wci_Vm_2_MFlag;

  // value method wci_Vm_3_mCmd
  output [2 : 0] wci_Vm_3_MCmd;

  // value method wci_Vm_3_mAddrSpace
  output wci_Vm_3_MAddrSpace;

  // value method wci_Vm_3_mByteEn
  output [3 : 0] wci_Vm_3_MByteEn;

  // value method wci_Vm_3_mAddr
  output [31 : 0] wci_Vm_3_MAddr;

  // value method wci_Vm_3_mData
  output [31 : 0] wci_Vm_3_MData;

  // action method wci_Vm_3_sResp
  input  [1 : 0] wci_Vm_3_SResp;

  // action method wci_Vm_3_sData
  input  [31 : 0] wci_Vm_3_SData;

  // action method wci_Vm_3_sThreadBusy
  input  wci_Vm_3_SThreadBusy;

  // action method wci_Vm_3_sFlag
  input  [2 : 0] wci_Vm_3_SFlag;

  // value method wci_Vm_3_mFlag
  output [1 : 0] wci_Vm_3_MFlag;

  // value method wci_Vm_4_mCmd
  output [2 : 0] wci_Vm_4_MCmd;

  // value method wci_Vm_4_mAddrSpace
  output wci_Vm_4_MAddrSpace;

  // value method wci_Vm_4_mByteEn
  output [3 : 0] wci_Vm_4_MByteEn;

  // value method wci_Vm_4_mAddr
  output [31 : 0] wci_Vm_4_MAddr;

  // value method wci_Vm_4_mData
  output [31 : 0] wci_Vm_4_MData;

  // action method wci_Vm_4_sResp
  input  [1 : 0] wci_Vm_4_SResp;

  // action method wci_Vm_4_sData
  input  [31 : 0] wci_Vm_4_SData;

  // action method wci_Vm_4_sThreadBusy
  input  wci_Vm_4_SThreadBusy;

  // action method wci_Vm_4_sFlag
  input  [2 : 0] wci_Vm_4_SFlag;

  // value method wci_Vm_4_mFlag
  output [1 : 0] wci_Vm_4_MFlag;

  // value method wci_Vm_5_mCmd
  output [2 : 0] wci_Vm_5_MCmd;

  // value method wci_Vm_5_mAddrSpace
  output wci_Vm_5_MAddrSpace;

  // value method wci_Vm_5_mByteEn
  output [3 : 0] wci_Vm_5_MByteEn;

  // value method wci_Vm_5_mAddr
  output [31 : 0] wci_Vm_5_MAddr;

  // value method wci_Vm_5_mData
  output [31 : 0] wci_Vm_5_MData;

  // action method wci_Vm_5_sResp
  input  [1 : 0] wci_Vm_5_SResp;

  // action method wci_Vm_5_sData
  input  [31 : 0] wci_Vm_5_SData;

  // action method wci_Vm_5_sThreadBusy
  input  wci_Vm_5_SThreadBusy;

  // action method wci_Vm_5_sFlag
  input  [2 : 0] wci_Vm_5_SFlag;

  // value method wci_Vm_5_mFlag
  output [1 : 0] wci_Vm_5_MFlag;

  // value method wci_Vm_6_mCmd
  output [2 : 0] wci_Vm_6_MCmd;

  // value method wci_Vm_6_mAddrSpace
  output wci_Vm_6_MAddrSpace;

  // value method wci_Vm_6_mByteEn
  output [3 : 0] wci_Vm_6_MByteEn;

  // value method wci_Vm_6_mAddr
  output [31 : 0] wci_Vm_6_MAddr;

  // value method wci_Vm_6_mData
  output [31 : 0] wci_Vm_6_MData;

  // action method wci_Vm_6_sResp
  input  [1 : 0] wci_Vm_6_SResp;

  // action method wci_Vm_6_sData
  input  [31 : 0] wci_Vm_6_SData;

  // action method wci_Vm_6_sThreadBusy
  input  wci_Vm_6_SThreadBusy;

  // action method wci_Vm_6_sFlag
  input  [2 : 0] wci_Vm_6_SFlag;

  // value method wci_Vm_6_mFlag
  output [1 : 0] wci_Vm_6_MFlag;

  // value method wci_Vm_7_mCmd
  output [2 : 0] wci_Vm_7_MCmd;

  // value method wci_Vm_7_mAddrSpace
  output wci_Vm_7_MAddrSpace;

  // value method wci_Vm_7_mByteEn
  output [3 : 0] wci_Vm_7_MByteEn;

  // value method wci_Vm_7_mAddr
  output [31 : 0] wci_Vm_7_MAddr;

  // value method wci_Vm_7_mData
  output [31 : 0] wci_Vm_7_MData;

  // action method wci_Vm_7_sResp
  input  [1 : 0] wci_Vm_7_SResp;

  // action method wci_Vm_7_sData
  input  [31 : 0] wci_Vm_7_SData;

  // action method wci_Vm_7_sThreadBusy
  input  wci_Vm_7_SThreadBusy;

  // action method wci_Vm_7_sFlag
  input  [2 : 0] wci_Vm_7_SFlag;

  // value method wci_Vm_7_mFlag
  output [1 : 0] wci_Vm_7_MFlag;

  // value method wci_Vm_8_mCmd
  output [2 : 0] wci_Vm_8_MCmd;

  // value method wci_Vm_8_mAddrSpace
  output wci_Vm_8_MAddrSpace;

  // value method wci_Vm_8_mByteEn
  output [3 : 0] wci_Vm_8_MByteEn;

  // value method wci_Vm_8_mAddr
  output [31 : 0] wci_Vm_8_MAddr;

  // value method wci_Vm_8_mData
  output [31 : 0] wci_Vm_8_MData;

  // action method wci_Vm_8_sResp
  input  [1 : 0] wci_Vm_8_SResp;

  // action method wci_Vm_8_sData
  input  [31 : 0] wci_Vm_8_SData;

  // action method wci_Vm_8_sThreadBusy
  input  wci_Vm_8_SThreadBusy;

  // action method wci_Vm_8_sFlag
  input  [2 : 0] wci_Vm_8_SFlag;

  // value method wci_Vm_8_mFlag
  output [1 : 0] wci_Vm_8_MFlag;

  // value method wci_Vm_9_mCmd
  output [2 : 0] wci_Vm_9_MCmd;

  // value method wci_Vm_9_mAddrSpace
  output wci_Vm_9_MAddrSpace;

  // value method wci_Vm_9_mByteEn
  output [3 : 0] wci_Vm_9_MByteEn;

  // value method wci_Vm_9_mAddr
  output [31 : 0] wci_Vm_9_MAddr;

  // value method wci_Vm_9_mData
  output [31 : 0] wci_Vm_9_MData;

  // action method wci_Vm_9_sResp
  input  [1 : 0] wci_Vm_9_SResp;

  // action method wci_Vm_9_sData
  input  [31 : 0] wci_Vm_9_SData;

  // action method wci_Vm_9_sThreadBusy
  input  wci_Vm_9_SThreadBusy;

  // action method wci_Vm_9_sFlag
  input  [2 : 0] wci_Vm_9_SFlag;

  // value method wci_Vm_9_mFlag
  output [1 : 0] wci_Vm_9_MFlag;

  // value method wci_Vm_10_mCmd
  output [2 : 0] wci_Vm_10_MCmd;

  // value method wci_Vm_10_mAddrSpace
  output wci_Vm_10_MAddrSpace;

  // value method wci_Vm_10_mByteEn
  output [3 : 0] wci_Vm_10_MByteEn;

  // value method wci_Vm_10_mAddr
  output [31 : 0] wci_Vm_10_MAddr;

  // value method wci_Vm_10_mData
  output [31 : 0] wci_Vm_10_MData;

  // action method wci_Vm_10_sResp
  input  [1 : 0] wci_Vm_10_SResp;

  // action method wci_Vm_10_sData
  input  [31 : 0] wci_Vm_10_SData;

  // action method wci_Vm_10_sThreadBusy
  input  wci_Vm_10_SThreadBusy;

  // action method wci_Vm_10_sFlag
  input  [2 : 0] wci_Vm_10_SFlag;

  // value method wci_Vm_10_mFlag
  output [1 : 0] wci_Vm_10_MFlag;

  // value method wci_Vm_11_mCmd
  output [2 : 0] wci_Vm_11_MCmd;

  // value method wci_Vm_11_mAddrSpace
  output wci_Vm_11_MAddrSpace;

  // value method wci_Vm_11_mByteEn
  output [3 : 0] wci_Vm_11_MByteEn;

  // value method wci_Vm_11_mAddr
  output [31 : 0] wci_Vm_11_MAddr;

  // value method wci_Vm_11_mData
  output [31 : 0] wci_Vm_11_MData;

  // action method wci_Vm_11_sResp
  input  [1 : 0] wci_Vm_11_SResp;

  // action method wci_Vm_11_sData
  input  [31 : 0] wci_Vm_11_SData;

  // action method wci_Vm_11_sThreadBusy
  input  wci_Vm_11_SThreadBusy;

  // action method wci_Vm_11_sFlag
  input  [2 : 0] wci_Vm_11_SFlag;

  // value method wci_Vm_11_mFlag
  output [1 : 0] wci_Vm_11_MFlag;

  // value method wci_Vm_12_mCmd
  output [2 : 0] wci_Vm_12_MCmd;

  // value method wci_Vm_12_mAddrSpace
  output wci_Vm_12_MAddrSpace;

  // value method wci_Vm_12_mByteEn
  output [3 : 0] wci_Vm_12_MByteEn;

  // value method wci_Vm_12_mAddr
  output [31 : 0] wci_Vm_12_MAddr;

  // value method wci_Vm_12_mData
  output [31 : 0] wci_Vm_12_MData;

  // action method wci_Vm_12_sResp
  input  [1 : 0] wci_Vm_12_SResp;

  // action method wci_Vm_12_sData
  input  [31 : 0] wci_Vm_12_SData;

  // action method wci_Vm_12_sThreadBusy
  input  wci_Vm_12_SThreadBusy;

  // action method wci_Vm_12_sFlag
  input  [2 : 0] wci_Vm_12_SFlag;

  // value method wci_Vm_12_mFlag
  output [1 : 0] wci_Vm_12_MFlag;

  // value method wci_Vm_13_mCmd
  output [2 : 0] wci_Vm_13_MCmd;

  // value method wci_Vm_13_mAddrSpace
  output wci_Vm_13_MAddrSpace;

  // value method wci_Vm_13_mByteEn
  output [3 : 0] wci_Vm_13_MByteEn;

  // value method wci_Vm_13_mAddr
  output [31 : 0] wci_Vm_13_MAddr;

  // value method wci_Vm_13_mData
  output [31 : 0] wci_Vm_13_MData;

  // action method wci_Vm_13_sResp
  input  [1 : 0] wci_Vm_13_SResp;

  // action method wci_Vm_13_sData
  input  [31 : 0] wci_Vm_13_SData;

  // action method wci_Vm_13_sThreadBusy
  input  wci_Vm_13_SThreadBusy;

  // action method wci_Vm_13_sFlag
  input  [2 : 0] wci_Vm_13_SFlag;

  // value method wci_Vm_13_mFlag
  output [1 : 0] wci_Vm_13_MFlag;

  // value method wci_Vm_14_mCmd
  output [2 : 0] wci_Vm_14_MCmd;

  // value method wci_Vm_14_mAddrSpace
  output wci_Vm_14_MAddrSpace;

  // value method wci_Vm_14_mByteEn
  output [3 : 0] wci_Vm_14_MByteEn;

  // value method wci_Vm_14_mAddr
  output [31 : 0] wci_Vm_14_MAddr;

  // value method wci_Vm_14_mData
  output [31 : 0] wci_Vm_14_MData;

  // action method wci_Vm_14_sResp
  input  [1 : 0] wci_Vm_14_SResp;

  // action method wci_Vm_14_sData
  input  [31 : 0] wci_Vm_14_SData;

  // action method wci_Vm_14_sThreadBusy
  input  wci_Vm_14_SThreadBusy;

  // action method wci_Vm_14_sFlag
  input  [2 : 0] wci_Vm_14_SFlag;

  // value method wci_Vm_14_mFlag
  output [1 : 0] wci_Vm_14_MFlag;

`ifdef not
  // value method cpNow
  output [63 : 0] cpNow;
  output RDY_cpNow;

  // action method gps_ppsSyncIn
  input  gps_ppsSyncIn_x;

  // value method gps_ppsSyncOut
  output gps_ppsSyncOut;

  // value method led
  output [1 : 0] led;

  // action method switch
  input  [2 : 0] switch_x;

  // action method uuid
  input  [511 : 0] uuid_arg;

  // Manually added metadata bram signals
  output       rom_en;
  output [9:0] rom_addr;
  input [31:0] rom_data;
`endif
  

  // output resets
  output RST_N_wci_Vm_0;
  output RST_N_wci_Vm_1;
  output RST_N_wci_Vm_2;
  output RST_N_wci_Vm_3;
  output RST_N_wci_Vm_4;
  output RST_N_wci_Vm_5;
  output RST_N_wci_Vm_6;
  output RST_N_wci_Vm_7;
  output RST_N_wci_Vm_8;
  output RST_N_wci_Vm_9;
  output RST_N_wci_Vm_10;
  output RST_N_wci_Vm_11;
  output RST_N_wci_Vm_12;
  output RST_N_wci_Vm_13;
  output RST_N_wci_Vm_14;

  // signals for module outputs
`ifdef not
  reg gps_ppsSyncOut;
  wire [63 : 0] cpNow;
`endif
  wire [39 : 0] server_response_get;
  wire [31 : 0] wci_Vm_0_MAddr,
		wci_Vm_0_MData,
		wci_Vm_10_MAddr,
		wci_Vm_10_MData,
		wci_Vm_11_MAddr,
		wci_Vm_11_MData,
		wci_Vm_12_MAddr,
		wci_Vm_12_MData,
		wci_Vm_13_MAddr,
		wci_Vm_13_MData,
		wci_Vm_14_MAddr,
		wci_Vm_14_MData,
		wci_Vm_1_MAddr,
		wci_Vm_1_MData,
		wci_Vm_2_MAddr,
		wci_Vm_2_MData,
		wci_Vm_3_MAddr,
		wci_Vm_3_MData,
		wci_Vm_4_MAddr,
		wci_Vm_4_MData,
		wci_Vm_5_MAddr,
		wci_Vm_5_MData,
		wci_Vm_6_MAddr,
		wci_Vm_6_MData,
		wci_Vm_7_MAddr,
		wci_Vm_7_MData,
		wci_Vm_8_MAddr,
		wci_Vm_8_MData,
		wci_Vm_9_MAddr,
		wci_Vm_9_MData;
  wire [3 : 0] wci_Vm_0_MByteEn,
	       wci_Vm_10_MByteEn,
	       wci_Vm_11_MByteEn,
	       wci_Vm_12_MByteEn,
	       wci_Vm_13_MByteEn,
	       wci_Vm_14_MByteEn,
	       wci_Vm_1_MByteEn,
	       wci_Vm_2_MByteEn,
	       wci_Vm_3_MByteEn,
	       wci_Vm_4_MByteEn,
	       wci_Vm_5_MByteEn,
	       wci_Vm_6_MByteEn,
	       wci_Vm_7_MByteEn,
	       wci_Vm_8_MByteEn,
	       wci_Vm_9_MByteEn;
  wire [2 : 0] wci_Vm_0_MCmd,
	       wci_Vm_10_MCmd,
	       wci_Vm_11_MCmd,
	       wci_Vm_12_MCmd,
	       wci_Vm_13_MCmd,
	       wci_Vm_14_MCmd,
	       wci_Vm_1_MCmd,
	       wci_Vm_2_MCmd,
	       wci_Vm_3_MCmd,
	       wci_Vm_4_MCmd,
	       wci_Vm_5_MCmd,
	       wci_Vm_6_MCmd,
	       wci_Vm_7_MCmd,
	       wci_Vm_8_MCmd,
	       wci_Vm_9_MCmd;
  wire [1 : 0] led,
	       wci_Vm_0_MFlag,
	       wci_Vm_10_MFlag,
	       wci_Vm_11_MFlag,
	       wci_Vm_12_MFlag,
	       wci_Vm_13_MFlag,
	       wci_Vm_14_MFlag,
	       wci_Vm_1_MFlag,
	       wci_Vm_2_MFlag,
	       wci_Vm_3_MFlag,
	       wci_Vm_4_MFlag,
	       wci_Vm_5_MFlag,
	       wci_Vm_6_MFlag,
	       wci_Vm_7_MFlag,
	       wci_Vm_8_MFlag,
	       wci_Vm_9_MFlag;
`ifdef not
  wire RDY_cpNow,
`else
  wire
`endif
       RDY_server_request_put,
       RDY_server_response_get,
       RST_N_wci_Vm_0,
       RST_N_wci_Vm_1,
       RST_N_wci_Vm_10,
       RST_N_wci_Vm_11,
       RST_N_wci_Vm_12,
       RST_N_wci_Vm_13,
       RST_N_wci_Vm_14,
       RST_N_wci_Vm_2,
       RST_N_wci_Vm_3,
       RST_N_wci_Vm_4,
       RST_N_wci_Vm_5,
       RST_N_wci_Vm_6,
       RST_N_wci_Vm_7,
       RST_N_wci_Vm_8,
       RST_N_wci_Vm_9,
       wci_Vm_0_MAddrSpace,
       wci_Vm_10_MAddrSpace,
       wci_Vm_11_MAddrSpace,
       wci_Vm_12_MAddrSpace,
       wci_Vm_13_MAddrSpace,
       wci_Vm_14_MAddrSpace,
       wci_Vm_1_MAddrSpace,
       wci_Vm_2_MAddrSpace,
       wci_Vm_3_MAddrSpace,
       wci_Vm_4_MAddrSpace,
       wci_Vm_5_MAddrSpace,
       wci_Vm_6_MAddrSpace,
       wci_Vm_7_MAddrSpace,
       wci_Vm_8_MAddrSpace,
       wci_Vm_9_MAddrSpace;

  // inlined wires
`ifdef not
  wire [511 : 0] uuidV$wget;
`endif
  wire [71 : 0] wci_reqF_10_x_wire$wget,
		wci_reqF_11_x_wire$wget,
		wci_reqF_12_x_wire$wget,
		wci_reqF_13_x_wire$wget,
		wci_reqF_14_x_wire$wget,
		wci_reqF_1_x_wire$wget,
		wci_reqF_2_x_wire$wget,
		wci_reqF_3_x_wire$wget,
		wci_reqF_4_x_wire$wget,
		wci_reqF_5_x_wire$wget,
		wci_reqF_6_x_wire$wget,
		wci_reqF_7_x_wire$wget,
		wci_reqF_8_x_wire$wget,
		wci_reqF_9_x_wire$wget,
		wci_reqF_x_wire$wget;
`ifdef not
  wire [63 : 0] devDNAV$wget, deviceDNA$wget;
  wire [49 : 0] timeServ_jamFracVal_1$wget;
`endif
  wire [33 : 0] wci_wciResponse$wget,
		wci_wciResponse_1$wget,
		wci_wciResponse_10$wget,
		wci_wciResponse_11$wget,
		wci_wciResponse_12$wget,
		wci_wciResponse_13$wget,
		wci_wciResponse_14$wget,
		wci_wciResponse_2$wget,
		wci_wciResponse_3$wget,
		wci_wciResponse_4$wget,
		wci_wciResponse_5$wget,
		wci_wciResponse_6$wget,
		wci_wciResponse_7$wget,
		wci_wciResponse_8$wget,
		wci_wciResponse_9$wget;
`ifdef not
  wire [31 : 0] rom_serverAdapter_outData_enqData$wget,
		rom_serverAdapter_outData_outData$wget,
`else
  wire [31 : 0]
`endif
		wci_Emv_respData_w$wget,
		wci_Emv_respData_w_1$wget,
		wci_Emv_respData_w_10$wget,
		wci_Emv_respData_w_11$wget,
		wci_Emv_respData_w_12$wget,
		wci_Emv_respData_w_13$wget,
		wci_Emv_respData_w_14$wget,
		wci_Emv_respData_w_2$wget,
		wci_Emv_respData_w_3$wget,
		wci_Emv_respData_w_4$wget,
		wci_Emv_respData_w_5$wget,
		wci_Emv_respData_w_6$wget,
		wci_Emv_respData_w_7$wget,
		wci_Emv_respData_w_8$wget,
		wci_Emv_respData_w_9$wget;
`ifdef not
  wire [2 : 0] rom_serverAdapter_cnt_1$wget,
	       rom_serverAdapter_cnt_2$wget,
	       rom_serverAdapter_cnt_3$wget;
  wire [1 : 0] rom_serverAdapter_s1_1$wget,
	       rom_serverAdapter_writeWithResp$wget,
`endif
  wire [1 : 0]	      
	       wci_Emv_resp_w$wget,
	       wci_Emv_resp_w_1$wget,
	       wci_Emv_resp_w_10$wget,
	       wci_Emv_resp_w_11$wget,
	       wci_Emv_resp_w_12$wget,
	       wci_Emv_resp_w_13$wget,
	       wci_Emv_resp_w_14$wget,
	       wci_Emv_resp_w_2$wget,
	       wci_Emv_resp_w_3$wget,
	       wci_Emv_resp_w_4$wget,
	       wci_Emv_resp_w_5$wget,
	       wci_Emv_resp_w_6$wget,
	       wci_Emv_resp_w_7$wget,
	       wci_Emv_resp_w_8$wget,
	       wci_Emv_resp_w_9$wget;
`ifdef not
  wire devDNAV$whas,
       deviceDNA$whas,
       dna_rdReg_1$wget,
       dna_rdReg_1$whas,
       dna_shftReg_1$wget,
       dna_shftReg_1$whas,
       rom_serverAdapter_cnt_1$whas,
       rom_serverAdapter_cnt_2$whas,
       rom_serverAdapter_cnt_3$whas,
       rom_serverAdapter_outData_deqCalled$whas,
       rom_serverAdapter_outData_enqData$whas,
       rom_serverAdapter_outData_outData$whas,
       rom_serverAdapter_s1_1$whas,
       rom_serverAdapter_writeWithResp$whas,
       timeServ_jamFracVal_1$whas,
       timeServ_jamFrac_1$wget,
       timeServ_jamFrac_1$whas,
       uuidV$whas,
`else
  wire 
`endif
       warmResetP_1$wget,
       warmResetP_1$whas,
       wci_Emv_respData_w$whas,
       wci_Emv_respData_w_1$whas,
       wci_Emv_respData_w_10$whas,
       wci_Emv_respData_w_11$whas,
       wci_Emv_respData_w_12$whas,
       wci_Emv_respData_w_13$whas,
       wci_Emv_respData_w_14$whas,
       wci_Emv_respData_w_2$whas,
       wci_Emv_respData_w_3$whas,
       wci_Emv_respData_w_4$whas,
       wci_Emv_respData_w_5$whas,
       wci_Emv_respData_w_6$whas,
       wci_Emv_respData_w_7$whas,
       wci_Emv_respData_w_8$whas,
       wci_Emv_respData_w_9$whas,
       wci_Emv_resp_w$whas,
       wci_Emv_resp_w_1$whas,
       wci_Emv_resp_w_10$whas,
       wci_Emv_resp_w_11$whas,
       wci_Emv_resp_w_12$whas,
       wci_Emv_resp_w_13$whas,
       wci_Emv_resp_w_14$whas,
       wci_Emv_resp_w_2$whas,
       wci_Emv_resp_w_3$whas,
       wci_Emv_resp_w_4$whas,
       wci_Emv_resp_w_5$whas,
       wci_Emv_resp_w_6$whas,
       wci_Emv_resp_w_7$whas,
       wci_Emv_resp_w_8$whas,
       wci_Emv_resp_w_9$whas,
       wci_reqF_10_dequeueing$whas,
       wci_reqF_10_enqueueing$whas,
       wci_reqF_10_x_wire$whas,
       wci_reqF_11_dequeueing$whas,
       wci_reqF_11_enqueueing$whas,
       wci_reqF_11_x_wire$whas,
       wci_reqF_12_dequeueing$whas,
       wci_reqF_12_enqueueing$whas,
       wci_reqF_12_x_wire$whas,
       wci_reqF_13_dequeueing$whas,
       wci_reqF_13_enqueueing$whas,
       wci_reqF_13_x_wire$whas,
       wci_reqF_14_dequeueing$whas,
       wci_reqF_14_enqueueing$whas,
       wci_reqF_14_x_wire$whas,
       wci_reqF_1_dequeueing$whas,
       wci_reqF_1_enqueueing$whas,
       wci_reqF_1_x_wire$whas,
       wci_reqF_2_dequeueing$whas,
       wci_reqF_2_enqueueing$whas,
       wci_reqF_2_x_wire$whas,
       wci_reqF_3_dequeueing$whas,
       wci_reqF_3_enqueueing$whas,
       wci_reqF_3_x_wire$whas,
       wci_reqF_4_dequeueing$whas,
       wci_reqF_4_enqueueing$whas,
       wci_reqF_4_x_wire$whas,
       wci_reqF_5_dequeueing$whas,
       wci_reqF_5_enqueueing$whas,
       wci_reqF_5_x_wire$whas,
       wci_reqF_6_dequeueing$whas,
       wci_reqF_6_enqueueing$whas,
       wci_reqF_6_x_wire$whas,
       wci_reqF_7_dequeueing$whas,
       wci_reqF_7_enqueueing$whas,
       wci_reqF_7_x_wire$whas,
       wci_reqF_8_dequeueing$whas,
       wci_reqF_8_enqueueing$whas,
       wci_reqF_8_x_wire$whas,
       wci_reqF_9_dequeueing$whas,
       wci_reqF_9_enqueueing$whas,
       wci_reqF_9_x_wire$whas,
       wci_reqF_dequeueing$whas,
       wci_reqF_enqueueing$whas,
       wci_reqF_x_wire$whas,
       wci_sThreadBusy_pw$whas,
       wci_sThreadBusy_pw_1$whas,
       wci_sThreadBusy_pw_10$whas,
       wci_sThreadBusy_pw_11$whas,
       wci_sThreadBusy_pw_12$whas,
       wci_sThreadBusy_pw_13$whas,
       wci_sThreadBusy_pw_14$whas,
       wci_sThreadBusy_pw_2$whas,
       wci_sThreadBusy_pw_3$whas,
       wci_sThreadBusy_pw_4$whas,
       wci_sThreadBusy_pw_5$whas,
       wci_sThreadBusy_pw_6$whas,
       wci_sThreadBusy_pw_7$whas,
       wci_sThreadBusy_pw_8$whas,
       wci_sThreadBusy_pw_9$whas,
       wci_sfCapClear_1$wget,
       wci_sfCapClear_1$whas,
       wci_sfCapClear_10_1$wget,
       wci_sfCapClear_10_1$whas,
       wci_sfCapClear_11_1$wget,
       wci_sfCapClear_11_1$whas,
       wci_sfCapClear_12_1$wget,
       wci_sfCapClear_12_1$whas,
       wci_sfCapClear_13_1$wget,
       wci_sfCapClear_13_1$whas,
       wci_sfCapClear_14_1$wget,
       wci_sfCapClear_14_1$whas,
       wci_sfCapClear_1_2$wget,
       wci_sfCapClear_1_2$whas,
       wci_sfCapClear_2_1$wget,
       wci_sfCapClear_2_1$whas,
       wci_sfCapClear_3_1$wget,
       wci_sfCapClear_3_1$whas,
       wci_sfCapClear_4_1$wget,
       wci_sfCapClear_4_1$whas,
       wci_sfCapClear_5_1$wget,
       wci_sfCapClear_5_1$whas,
       wci_sfCapClear_6_1$wget,
       wci_sfCapClear_6_1$whas,
       wci_sfCapClear_7_1$wget,
       wci_sfCapClear_7_1$whas,
       wci_sfCapClear_8_1$wget,
       wci_sfCapClear_8_1$whas,
       wci_sfCapClear_9_1$wget,
       wci_sfCapClear_9_1$whas,
       wci_sfCapSet_1$wget,
       wci_sfCapSet_1$whas,
       wci_sfCapSet_10_1$wget,
       wci_sfCapSet_10_1$whas,
       wci_sfCapSet_11_1$wget,
       wci_sfCapSet_11_1$whas,
       wci_sfCapSet_12_1$wget,
       wci_sfCapSet_12_1$whas,
       wci_sfCapSet_13_1$wget,
       wci_sfCapSet_13_1$whas,
       wci_sfCapSet_14_1$wget,
       wci_sfCapSet_14_1$whas,
       wci_sfCapSet_1_2$wget,
       wci_sfCapSet_1_2$whas,
       wci_sfCapSet_2_1$wget,
       wci_sfCapSet_2_1$whas,
       wci_sfCapSet_3_1$wget,
       wci_sfCapSet_3_1$whas,
       wci_sfCapSet_4_1$wget,
       wci_sfCapSet_4_1$whas,
       wci_sfCapSet_5_1$wget,
       wci_sfCapSet_5_1$whas,
       wci_sfCapSet_6_1$wget,
       wci_sfCapSet_6_1$whas,
       wci_sfCapSet_7_1$wget,
       wci_sfCapSet_7_1$whas,
       wci_sfCapSet_8_1$wget,
       wci_sfCapSet_8_1$whas,
       wci_sfCapSet_9_1$wget,
       wci_sfCapSet_9_1$whas,
       wci_wciResponse$whas,
       wci_wciResponse_1$whas,
       wci_wciResponse_10$whas,
       wci_wciResponse_11$whas,
       wci_wciResponse_12$whas,
       wci_wciResponse_13$whas,
       wci_wciResponse_14$whas,
       wci_wciResponse_2$whas,
       wci_wciResponse_3$whas,
       wci_wciResponse_4$whas,
       wci_wciResponse_5$whas,
       wci_wciResponse_6$whas,
       wci_wciResponse_7$whas,
       wci_wciResponse_8$whas,
       wci_wciResponse_9$whas;

  // register cpControl
  reg [31 : 0] cpControl;
  wire [31 : 0] cpControl$D_IN;
  wire cpControl$EN;

  // register cpReq
  reg [64 : 0] cpReq;
  reg [64 : 0] cpReq$D_IN;
  wire cpReq$EN;

`ifdef not
  // register deltaTime
  reg [63 : 0] deltaTime;
  wire [63 : 0] deltaTime$D_IN;
  wire deltaTime$EN;
`endif

  // register dispatched
  reg dispatched;
  reg dispatched$D_IN;
  wire dispatched$EN;

`ifdef not
  // register dna_cnt
  reg [6 : 0] dna_cnt;
  wire [6 : 0] dna_cnt$D_IN;
  wire dna_cnt$EN;

  // register dna_rdReg
  reg dna_rdReg;
  wire dna_rdReg$D_IN, dna_rdReg$EN;

  // register dna_shftReg
  reg dna_shftReg;
  wire dna_shftReg$D_IN, dna_shftReg$EN;

  // register dna_sr
  reg [56 : 0] dna_sr;
  wire [56 : 0] dna_sr$D_IN;
  wire dna_sr$EN;
`endif

  // register readCntReg
  reg [31 : 0] readCntReg;
  wire [31 : 0] readCntReg$D_IN;
  wire readCntReg$EN;

  // register rogueTLP
  reg [3 : 0] rogueTLP;
  wire [3 : 0] rogueTLP$D_IN;
  wire rogueTLP$EN;

`ifdef not
  // register rom_serverAdapter_cnt
  reg [2 : 0] rom_serverAdapter_cnt;
  wire [2 : 0] rom_serverAdapter_cnt$D_IN;
  wire rom_serverAdapter_cnt$EN;

  // register rom_serverAdapter_s1
  reg [1 : 0] rom_serverAdapter_s1;
  wire [1 : 0] rom_serverAdapter_s1$D_IN;
  wire rom_serverAdapter_s1$EN;
`endif

  // register scratch20
  reg [31 : 0] scratch20;
  wire [31 : 0] scratch20$D_IN;
  wire scratch20$EN;

  // register scratch24
  reg [31 : 0] scratch24;
  wire [31 : 0] scratch24$D_IN;
  wire scratch24$EN;

  // register seqTag
  reg [7 : 0] seqTag;
  wire [7 : 0] seqTag$D_IN;
  wire seqTag$EN;

`ifdef not
  // register switch_d
  reg [2 : 0] switch_d;
  wire [2 : 0] switch_d$D_IN;
  wire switch_d$EN;
`endif

  // register td
  reg [31 : 0] td;
  wire [31 : 0] td$D_IN;
  wire td$EN;

`ifdef not
  // register timeServ_delSec
  reg [1 : 0] timeServ_delSec;
  wire [1 : 0] timeServ_delSec$D_IN;
  wire timeServ_delSec$EN;

  // register timeServ_delSecond
  reg [49 : 0] timeServ_delSecond;
  wire [49 : 0] timeServ_delSecond$D_IN;
  wire timeServ_delSecond$EN;

  // register timeServ_fracInc
  reg [49 : 0] timeServ_fracInc;
  wire [49 : 0] timeServ_fracInc$D_IN;
  wire timeServ_fracInc$EN;

  // register timeServ_fracSeconds
  reg [49 : 0] timeServ_fracSeconds;
  wire [49 : 0] timeServ_fracSeconds$D_IN;
  wire timeServ_fracSeconds$EN;

  // register timeServ_gpsInSticky
  reg timeServ_gpsInSticky;
  wire timeServ_gpsInSticky$D_IN, timeServ_gpsInSticky$EN;

  // register timeServ_jamFrac
  reg timeServ_jamFrac;
  wire timeServ_jamFrac$D_IN, timeServ_jamFrac$EN;

  // register timeServ_jamFracVal
  reg [49 : 0] timeServ_jamFracVal;
  wire [49 : 0] timeServ_jamFracVal$D_IN;
  wire timeServ_jamFracVal$EN;

  // register timeServ_lastSecond
  reg [49 : 0] timeServ_lastSecond;
  wire [49 : 0] timeServ_lastSecond$D_IN;
  wire timeServ_lastSecond$EN;

  // register timeServ_now
  reg [63 : 0] timeServ_now;
  wire [63 : 0] timeServ_now$D_IN;
  wire timeServ_now$EN;

  // register timeServ_ppsDrive
  reg timeServ_ppsDrive;
  wire timeServ_ppsDrive$D_IN, timeServ_ppsDrive$EN;

  // register timeServ_ppsEdgeCount
  reg [7 : 0] timeServ_ppsEdgeCount;
  wire [7 : 0] timeServ_ppsEdgeCount$D_IN;
  wire timeServ_ppsEdgeCount$EN;

  // register timeServ_ppsExtCapture
  reg timeServ_ppsExtCapture;
  wire timeServ_ppsExtCapture$D_IN, timeServ_ppsExtCapture$EN;

  // register timeServ_ppsExtSyncD
  reg timeServ_ppsExtSyncD;
  wire timeServ_ppsExtSyncD$D_IN, timeServ_ppsExtSyncD$EN;

  // register timeServ_ppsExtSync_d1
  reg timeServ_ppsExtSync_d1;
  wire timeServ_ppsExtSync_d1$D_IN, timeServ_ppsExtSync_d1$EN;

  // register timeServ_ppsExtSync_d2
  reg timeServ_ppsExtSync_d2;
  wire timeServ_ppsExtSync_d2$D_IN, timeServ_ppsExtSync_d2$EN;

  // register timeServ_ppsInSticky
  reg timeServ_ppsInSticky;
  wire timeServ_ppsInSticky$D_IN, timeServ_ppsInSticky$EN;

  // register timeServ_ppsLost
  reg timeServ_ppsLost;
  wire timeServ_ppsLost$D_IN, timeServ_ppsLost$EN;

  // register timeServ_ppsLostSticky
  reg timeServ_ppsLostSticky;
  wire timeServ_ppsLostSticky$D_IN, timeServ_ppsLostSticky$EN;

  // register timeServ_ppsOK
  reg timeServ_ppsOK;
  wire timeServ_ppsOK$D_IN, timeServ_ppsOK$EN;

  // register timeServ_refFreeCount
  reg [27 : 0] timeServ_refFreeCount;
  wire [27 : 0] timeServ_refFreeCount$D_IN;
  wire timeServ_refFreeCount$EN;

  // register timeServ_refFreeSamp
  reg [27 : 0] timeServ_refFreeSamp;
  wire [27 : 0] timeServ_refFreeSamp$D_IN;
  wire timeServ_refFreeSamp$EN;

  // register timeServ_refFreeSpan
  reg [27 : 0] timeServ_refFreeSpan;
  wire [27 : 0] timeServ_refFreeSpan$D_IN;
  wire timeServ_refFreeSpan$EN;

  // register timeServ_refFromRise
  reg [27 : 0] timeServ_refFromRise;
  wire [27 : 0] timeServ_refFromRise$D_IN;
  wire timeServ_refFromRise$EN;

  // register timeServ_refPerCount
  reg [27 : 0] timeServ_refPerCount;
  wire [27 : 0] timeServ_refPerCount$D_IN;
  wire timeServ_refPerCount$EN;

  // register timeServ_refSecCount
  reg [31 : 0] timeServ_refSecCount;
  wire [31 : 0] timeServ_refSecCount$D_IN;
  wire timeServ_refSecCount$EN;

  // register timeServ_rplTimeControl
  reg [4 : 0] timeServ_rplTimeControl;
  wire [4 : 0] timeServ_rplTimeControl$D_IN;
  wire timeServ_rplTimeControl$EN;

  // register timeServ_timeSetSticky
  reg timeServ_timeSetSticky;
  wire timeServ_timeSetSticky$D_IN, timeServ_timeSetSticky$EN;

  // register timeServ_xo2
  reg timeServ_xo2;
  wire timeServ_xo2$D_IN, timeServ_xo2$EN;
`endif

  // register warmResetP
  reg warmResetP;
  wire warmResetP$D_IN, warmResetP$EN;

  // register wci_busy
  reg wci_busy;
  wire wci_busy$D_IN, wci_busy$EN;

  // register wci_busy_1
  reg wci_busy_1;
  wire wci_busy_1$D_IN, wci_busy_1$EN;

  // register wci_busy_10
  reg wci_busy_10;
  wire wci_busy_10$D_IN, wci_busy_10$EN;

  // register wci_busy_11
  reg wci_busy_11;
  wire wci_busy_11$D_IN, wci_busy_11$EN;

  // register wci_busy_12
  reg wci_busy_12;
  wire wci_busy_12$D_IN, wci_busy_12$EN;

  // register wci_busy_13
  reg wci_busy_13;
  wire wci_busy_13$D_IN, wci_busy_13$EN;

  // register wci_busy_14
  reg wci_busy_14;
  wire wci_busy_14$D_IN, wci_busy_14$EN;

  // register wci_busy_2
  reg wci_busy_2;
  wire wci_busy_2$D_IN, wci_busy_2$EN;

  // register wci_busy_3
  reg wci_busy_3;
  wire wci_busy_3$D_IN, wci_busy_3$EN;

  // register wci_busy_4
  reg wci_busy_4;
  wire wci_busy_4$D_IN, wci_busy_4$EN;

  // register wci_busy_5
  reg wci_busy_5;
  wire wci_busy_5$D_IN, wci_busy_5$EN;

  // register wci_busy_6
  reg wci_busy_6;
  wire wci_busy_6$D_IN, wci_busy_6$EN;

  // register wci_busy_7
  reg wci_busy_7;
  wire wci_busy_7$D_IN, wci_busy_7$EN;

  // register wci_busy_8
  reg wci_busy_8;
  wire wci_busy_8$D_IN, wci_busy_8$EN;

  // register wci_busy_9
  reg wci_busy_9;
  wire wci_busy_9$D_IN, wci_busy_9$EN;

  // register wci_lastConfigAddr
  reg [32 : 0] wci_lastConfigAddr;
  wire [32 : 0] wci_lastConfigAddr$D_IN;
  wire wci_lastConfigAddr$EN;

  // register wci_lastConfigAddr_1
  reg [32 : 0] wci_lastConfigAddr_1;
  wire [32 : 0] wci_lastConfigAddr_1$D_IN;
  wire wci_lastConfigAddr_1$EN;

  // register wci_lastConfigAddr_10
  reg [32 : 0] wci_lastConfigAddr_10;
  wire [32 : 0] wci_lastConfigAddr_10$D_IN;
  wire wci_lastConfigAddr_10$EN;

  // register wci_lastConfigAddr_11
  reg [32 : 0] wci_lastConfigAddr_11;
  wire [32 : 0] wci_lastConfigAddr_11$D_IN;
  wire wci_lastConfigAddr_11$EN;

  // register wci_lastConfigAddr_12
  reg [32 : 0] wci_lastConfigAddr_12;
  wire [32 : 0] wci_lastConfigAddr_12$D_IN;
  wire wci_lastConfigAddr_12$EN;

  // register wci_lastConfigAddr_13
  reg [32 : 0] wci_lastConfigAddr_13;
  wire [32 : 0] wci_lastConfigAddr_13$D_IN;
  wire wci_lastConfigAddr_13$EN;

  // register wci_lastConfigAddr_14
  reg [32 : 0] wci_lastConfigAddr_14;
  wire [32 : 0] wci_lastConfigAddr_14$D_IN;
  wire wci_lastConfigAddr_14$EN;

  // register wci_lastConfigAddr_2
  reg [32 : 0] wci_lastConfigAddr_2;
  wire [32 : 0] wci_lastConfigAddr_2$D_IN;
  wire wci_lastConfigAddr_2$EN;

  // register wci_lastConfigAddr_3
  reg [32 : 0] wci_lastConfigAddr_3;
  wire [32 : 0] wci_lastConfigAddr_3$D_IN;
  wire wci_lastConfigAddr_3$EN;

  // register wci_lastConfigAddr_4
  reg [32 : 0] wci_lastConfigAddr_4;
  wire [32 : 0] wci_lastConfigAddr_4$D_IN;
  wire wci_lastConfigAddr_4$EN;

  // register wci_lastConfigAddr_5
  reg [32 : 0] wci_lastConfigAddr_5;
  wire [32 : 0] wci_lastConfigAddr_5$D_IN;
  wire wci_lastConfigAddr_5$EN;

  // register wci_lastConfigAddr_6
  reg [32 : 0] wci_lastConfigAddr_6;
  wire [32 : 0] wci_lastConfigAddr_6$D_IN;
  wire wci_lastConfigAddr_6$EN;

  // register wci_lastConfigAddr_7
  reg [32 : 0] wci_lastConfigAddr_7;
  wire [32 : 0] wci_lastConfigAddr_7$D_IN;
  wire wci_lastConfigAddr_7$EN;

  // register wci_lastConfigAddr_8
  reg [32 : 0] wci_lastConfigAddr_8;
  wire [32 : 0] wci_lastConfigAddr_8$D_IN;
  wire wci_lastConfigAddr_8$EN;

  // register wci_lastConfigAddr_9
  reg [32 : 0] wci_lastConfigAddr_9;
  wire [32 : 0] wci_lastConfigAddr_9$D_IN;
  wire wci_lastConfigAddr_9$EN;

  // register wci_lastConfigBE
  reg [4 : 0] wci_lastConfigBE;
  wire [4 : 0] wci_lastConfigBE$D_IN;
  wire wci_lastConfigBE$EN;

  // register wci_lastConfigBE_1
  reg [4 : 0] wci_lastConfigBE_1;
  wire [4 : 0] wci_lastConfigBE_1$D_IN;
  wire wci_lastConfigBE_1$EN;

  // register wci_lastConfigBE_10
  reg [4 : 0] wci_lastConfigBE_10;
  wire [4 : 0] wci_lastConfigBE_10$D_IN;
  wire wci_lastConfigBE_10$EN;

  // register wci_lastConfigBE_11
  reg [4 : 0] wci_lastConfigBE_11;
  wire [4 : 0] wci_lastConfigBE_11$D_IN;
  wire wci_lastConfigBE_11$EN;

  // register wci_lastConfigBE_12
  reg [4 : 0] wci_lastConfigBE_12;
  wire [4 : 0] wci_lastConfigBE_12$D_IN;
  wire wci_lastConfigBE_12$EN;

  // register wci_lastConfigBE_13
  reg [4 : 0] wci_lastConfigBE_13;
  wire [4 : 0] wci_lastConfigBE_13$D_IN;
  wire wci_lastConfigBE_13$EN;

  // register wci_lastConfigBE_14
  reg [4 : 0] wci_lastConfigBE_14;
  wire [4 : 0] wci_lastConfigBE_14$D_IN;
  wire wci_lastConfigBE_14$EN;

  // register wci_lastConfigBE_2
  reg [4 : 0] wci_lastConfigBE_2;
  wire [4 : 0] wci_lastConfigBE_2$D_IN;
  wire wci_lastConfigBE_2$EN;

  // register wci_lastConfigBE_3
  reg [4 : 0] wci_lastConfigBE_3;
  wire [4 : 0] wci_lastConfigBE_3$D_IN;
  wire wci_lastConfigBE_3$EN;

  // register wci_lastConfigBE_4
  reg [4 : 0] wci_lastConfigBE_4;
  wire [4 : 0] wci_lastConfigBE_4$D_IN;
  wire wci_lastConfigBE_4$EN;

  // register wci_lastConfigBE_5
  reg [4 : 0] wci_lastConfigBE_5;
  wire [4 : 0] wci_lastConfigBE_5$D_IN;
  wire wci_lastConfigBE_5$EN;

  // register wci_lastConfigBE_6
  reg [4 : 0] wci_lastConfigBE_6;
  wire [4 : 0] wci_lastConfigBE_6$D_IN;
  wire wci_lastConfigBE_6$EN;

  // register wci_lastConfigBE_7
  reg [4 : 0] wci_lastConfigBE_7;
  wire [4 : 0] wci_lastConfigBE_7$D_IN;
  wire wci_lastConfigBE_7$EN;

  // register wci_lastConfigBE_8
  reg [4 : 0] wci_lastConfigBE_8;
  wire [4 : 0] wci_lastConfigBE_8$D_IN;
  wire wci_lastConfigBE_8$EN;

  // register wci_lastConfigBE_9
  reg [4 : 0] wci_lastConfigBE_9;
  wire [4 : 0] wci_lastConfigBE_9$D_IN;
  wire wci_lastConfigBE_9$EN;

  // register wci_lastControlOp
  reg [3 : 0] wci_lastControlOp;
  wire [3 : 0] wci_lastControlOp$D_IN;
  wire wci_lastControlOp$EN;

  // register wci_lastControlOp_1
  reg [3 : 0] wci_lastControlOp_1;
  wire [3 : 0] wci_lastControlOp_1$D_IN;
  wire wci_lastControlOp_1$EN;

  // register wci_lastControlOp_10
  reg [3 : 0] wci_lastControlOp_10;
  wire [3 : 0] wci_lastControlOp_10$D_IN;
  wire wci_lastControlOp_10$EN;

  // register wci_lastControlOp_11
  reg [3 : 0] wci_lastControlOp_11;
  wire [3 : 0] wci_lastControlOp_11$D_IN;
  wire wci_lastControlOp_11$EN;

  // register wci_lastControlOp_12
  reg [3 : 0] wci_lastControlOp_12;
  wire [3 : 0] wci_lastControlOp_12$D_IN;
  wire wci_lastControlOp_12$EN;

  // register wci_lastControlOp_13
  reg [3 : 0] wci_lastControlOp_13;
  wire [3 : 0] wci_lastControlOp_13$D_IN;
  wire wci_lastControlOp_13$EN;

  // register wci_lastControlOp_14
  reg [3 : 0] wci_lastControlOp_14;
  wire [3 : 0] wci_lastControlOp_14$D_IN;
  wire wci_lastControlOp_14$EN;

  // register wci_lastControlOp_2
  reg [3 : 0] wci_lastControlOp_2;
  wire [3 : 0] wci_lastControlOp_2$D_IN;
  wire wci_lastControlOp_2$EN;

  // register wci_lastControlOp_3
  reg [3 : 0] wci_lastControlOp_3;
  wire [3 : 0] wci_lastControlOp_3$D_IN;
  wire wci_lastControlOp_3$EN;

  // register wci_lastControlOp_4
  reg [3 : 0] wci_lastControlOp_4;
  wire [3 : 0] wci_lastControlOp_4$D_IN;
  wire wci_lastControlOp_4$EN;

  // register wci_lastControlOp_5
  reg [3 : 0] wci_lastControlOp_5;
  wire [3 : 0] wci_lastControlOp_5$D_IN;
  wire wci_lastControlOp_5$EN;

  // register wci_lastControlOp_6
  reg [3 : 0] wci_lastControlOp_6;
  wire [3 : 0] wci_lastControlOp_6$D_IN;
  wire wci_lastControlOp_6$EN;

  // register wci_lastControlOp_7
  reg [3 : 0] wci_lastControlOp_7;
  wire [3 : 0] wci_lastControlOp_7$D_IN;
  wire wci_lastControlOp_7$EN;

  // register wci_lastControlOp_8
  reg [3 : 0] wci_lastControlOp_8;
  wire [3 : 0] wci_lastControlOp_8$D_IN;
  wire wci_lastControlOp_8$EN;

  // register wci_lastControlOp_9
  reg [3 : 0] wci_lastControlOp_9;
  wire [3 : 0] wci_lastControlOp_9$D_IN;
  wire wci_lastControlOp_9$EN;

  // register wci_lastOpWrite
  reg [1 : 0] wci_lastOpWrite;
  wire [1 : 0] wci_lastOpWrite$D_IN;
  wire wci_lastOpWrite$EN;

  // register wci_lastOpWrite_1
  reg [1 : 0] wci_lastOpWrite_1;
  wire [1 : 0] wci_lastOpWrite_1$D_IN;
  wire wci_lastOpWrite_1$EN;

  // register wci_lastOpWrite_10
  reg [1 : 0] wci_lastOpWrite_10;
  wire [1 : 0] wci_lastOpWrite_10$D_IN;
  wire wci_lastOpWrite_10$EN;

  // register wci_lastOpWrite_11
  reg [1 : 0] wci_lastOpWrite_11;
  wire [1 : 0] wci_lastOpWrite_11$D_IN;
  wire wci_lastOpWrite_11$EN;

  // register wci_lastOpWrite_12
  reg [1 : 0] wci_lastOpWrite_12;
  wire [1 : 0] wci_lastOpWrite_12$D_IN;
  wire wci_lastOpWrite_12$EN;

  // register wci_lastOpWrite_13
  reg [1 : 0] wci_lastOpWrite_13;
  wire [1 : 0] wci_lastOpWrite_13$D_IN;
  wire wci_lastOpWrite_13$EN;

  // register wci_lastOpWrite_14
  reg [1 : 0] wci_lastOpWrite_14;
  wire [1 : 0] wci_lastOpWrite_14$D_IN;
  wire wci_lastOpWrite_14$EN;

  // register wci_lastOpWrite_2
  reg [1 : 0] wci_lastOpWrite_2;
  wire [1 : 0] wci_lastOpWrite_2$D_IN;
  wire wci_lastOpWrite_2$EN;

  // register wci_lastOpWrite_3
  reg [1 : 0] wci_lastOpWrite_3;
  wire [1 : 0] wci_lastOpWrite_3$D_IN;
  wire wci_lastOpWrite_3$EN;

  // register wci_lastOpWrite_4
  reg [1 : 0] wci_lastOpWrite_4;
  wire [1 : 0] wci_lastOpWrite_4$D_IN;
  wire wci_lastOpWrite_4$EN;

  // register wci_lastOpWrite_5
  reg [1 : 0] wci_lastOpWrite_5;
  wire [1 : 0] wci_lastOpWrite_5$D_IN;
  wire wci_lastOpWrite_5$EN;

  // register wci_lastOpWrite_6
  reg [1 : 0] wci_lastOpWrite_6;
  wire [1 : 0] wci_lastOpWrite_6$D_IN;
  wire wci_lastOpWrite_6$EN;

  // register wci_lastOpWrite_7
  reg [1 : 0] wci_lastOpWrite_7;
  wire [1 : 0] wci_lastOpWrite_7$D_IN;
  wire wci_lastOpWrite_7$EN;

  // register wci_lastOpWrite_8
  reg [1 : 0] wci_lastOpWrite_8;
  wire [1 : 0] wci_lastOpWrite_8$D_IN;
  wire wci_lastOpWrite_8$EN;

  // register wci_lastOpWrite_9
  reg [1 : 0] wci_lastOpWrite_9;
  wire [1 : 0] wci_lastOpWrite_9$D_IN;
  wire wci_lastOpWrite_9$EN;

  // register wci_mFlagReg
  reg [1 : 0] wci_mFlagReg;
  wire [1 : 0] wci_mFlagReg$D_IN;
  wire wci_mFlagReg$EN;

  // register wci_mFlagReg_1
  reg [1 : 0] wci_mFlagReg_1;
  wire [1 : 0] wci_mFlagReg_1$D_IN;
  wire wci_mFlagReg_1$EN;

  // register wci_mFlagReg_10
  reg [1 : 0] wci_mFlagReg_10;
  wire [1 : 0] wci_mFlagReg_10$D_IN;
  wire wci_mFlagReg_10$EN;

  // register wci_mFlagReg_11
  reg [1 : 0] wci_mFlagReg_11;
  wire [1 : 0] wci_mFlagReg_11$D_IN;
  wire wci_mFlagReg_11$EN;

  // register wci_mFlagReg_12
  reg [1 : 0] wci_mFlagReg_12;
  wire [1 : 0] wci_mFlagReg_12$D_IN;
  wire wci_mFlagReg_12$EN;

  // register wci_mFlagReg_13
  reg [1 : 0] wci_mFlagReg_13;
  wire [1 : 0] wci_mFlagReg_13$D_IN;
  wire wci_mFlagReg_13$EN;

  // register wci_mFlagReg_14
  reg [1 : 0] wci_mFlagReg_14;
  wire [1 : 0] wci_mFlagReg_14$D_IN;
  wire wci_mFlagReg_14$EN;

  // register wci_mFlagReg_2
  reg [1 : 0] wci_mFlagReg_2;
  wire [1 : 0] wci_mFlagReg_2$D_IN;
  wire wci_mFlagReg_2$EN;

  // register wci_mFlagReg_3
  reg [1 : 0] wci_mFlagReg_3;
  wire [1 : 0] wci_mFlagReg_3$D_IN;
  wire wci_mFlagReg_3$EN;

  // register wci_mFlagReg_4
  reg [1 : 0] wci_mFlagReg_4;
  wire [1 : 0] wci_mFlagReg_4$D_IN;
  wire wci_mFlagReg_4$EN;

  // register wci_mFlagReg_5
  reg [1 : 0] wci_mFlagReg_5;
  wire [1 : 0] wci_mFlagReg_5$D_IN;
  wire wci_mFlagReg_5$EN;

  // register wci_mFlagReg_6
  reg [1 : 0] wci_mFlagReg_6;
  wire [1 : 0] wci_mFlagReg_6$D_IN;
  wire wci_mFlagReg_6$EN;

  // register wci_mFlagReg_7
  reg [1 : 0] wci_mFlagReg_7;
  wire [1 : 0] wci_mFlagReg_7$D_IN;
  wire wci_mFlagReg_7$EN;

  // register wci_mFlagReg_8
  reg [1 : 0] wci_mFlagReg_8;
  wire [1 : 0] wci_mFlagReg_8$D_IN;
  wire wci_mFlagReg_8$EN;

  // register wci_mFlagReg_9
  reg [1 : 0] wci_mFlagReg_9;
  wire [1 : 0] wci_mFlagReg_9$D_IN;
  wire wci_mFlagReg_9$EN;

  // register wci_pageWindow
  reg [11 : 0] wci_pageWindow;
  wire [11 : 0] wci_pageWindow$D_IN;
  wire wci_pageWindow$EN;

  // register wci_pageWindow_1
  reg [11 : 0] wci_pageWindow_1;
  wire [11 : 0] wci_pageWindow_1$D_IN;
  wire wci_pageWindow_1$EN;

  // register wci_pageWindow_10
  reg [11 : 0] wci_pageWindow_10;
  wire [11 : 0] wci_pageWindow_10$D_IN;
  wire wci_pageWindow_10$EN;

  // register wci_pageWindow_11
  reg [11 : 0] wci_pageWindow_11;
  wire [11 : 0] wci_pageWindow_11$D_IN;
  wire wci_pageWindow_11$EN;

  // register wci_pageWindow_12
  reg [11 : 0] wci_pageWindow_12;
  wire [11 : 0] wci_pageWindow_12$D_IN;
  wire wci_pageWindow_12$EN;

  // register wci_pageWindow_13
  reg [11 : 0] wci_pageWindow_13;
  wire [11 : 0] wci_pageWindow_13$D_IN;
  wire wci_pageWindow_13$EN;

  // register wci_pageWindow_14
  reg [11 : 0] wci_pageWindow_14;
  wire [11 : 0] wci_pageWindow_14$D_IN;
  wire wci_pageWindow_14$EN;

  // register wci_pageWindow_2
  reg [11 : 0] wci_pageWindow_2;
  wire [11 : 0] wci_pageWindow_2$D_IN;
  wire wci_pageWindow_2$EN;

  // register wci_pageWindow_3
  reg [11 : 0] wci_pageWindow_3;
  wire [11 : 0] wci_pageWindow_3$D_IN;
  wire wci_pageWindow_3$EN;

  // register wci_pageWindow_4
  reg [11 : 0] wci_pageWindow_4;
  wire [11 : 0] wci_pageWindow_4$D_IN;
  wire wci_pageWindow_4$EN;

  // register wci_pageWindow_5
  reg [11 : 0] wci_pageWindow_5;
  wire [11 : 0] wci_pageWindow_5$D_IN;
  wire wci_pageWindow_5$EN;

  // register wci_pageWindow_6
  reg [11 : 0] wci_pageWindow_6;
  wire [11 : 0] wci_pageWindow_6$D_IN;
  wire wci_pageWindow_6$EN;

  // register wci_pageWindow_7
  reg [11 : 0] wci_pageWindow_7;
  wire [11 : 0] wci_pageWindow_7$D_IN;
  wire wci_pageWindow_7$EN;

  // register wci_pageWindow_8
  reg [11 : 0] wci_pageWindow_8;
  wire [11 : 0] wci_pageWindow_8$D_IN;
  wire wci_pageWindow_8$EN;

  // register wci_pageWindow_9
  reg [11 : 0] wci_pageWindow_9;
  wire [11 : 0] wci_pageWindow_9$D_IN;
  wire wci_pageWindow_9$EN;

  // register wci_reqERR
  reg [2 : 0] wci_reqERR;
  wire [2 : 0] wci_reqERR$D_IN;
  wire wci_reqERR$EN;

  // register wci_reqERR_1
  reg [2 : 0] wci_reqERR_1;
  wire [2 : 0] wci_reqERR_1$D_IN;
  wire wci_reqERR_1$EN;

  // register wci_reqERR_10
  reg [2 : 0] wci_reqERR_10;
  wire [2 : 0] wci_reqERR_10$D_IN;
  wire wci_reqERR_10$EN;

  // register wci_reqERR_11
  reg [2 : 0] wci_reqERR_11;
  wire [2 : 0] wci_reqERR_11$D_IN;
  wire wci_reqERR_11$EN;

  // register wci_reqERR_12
  reg [2 : 0] wci_reqERR_12;
  wire [2 : 0] wci_reqERR_12$D_IN;
  wire wci_reqERR_12$EN;

  // register wci_reqERR_13
  reg [2 : 0] wci_reqERR_13;
  wire [2 : 0] wci_reqERR_13$D_IN;
  wire wci_reqERR_13$EN;

  // register wci_reqERR_14
  reg [2 : 0] wci_reqERR_14;
  wire [2 : 0] wci_reqERR_14$D_IN;
  wire wci_reqERR_14$EN;

  // register wci_reqERR_2
  reg [2 : 0] wci_reqERR_2;
  wire [2 : 0] wci_reqERR_2$D_IN;
  wire wci_reqERR_2$EN;

  // register wci_reqERR_3
  reg [2 : 0] wci_reqERR_3;
  wire [2 : 0] wci_reqERR_3$D_IN;
  wire wci_reqERR_3$EN;

  // register wci_reqERR_4
  reg [2 : 0] wci_reqERR_4;
  wire [2 : 0] wci_reqERR_4$D_IN;
  wire wci_reqERR_4$EN;

  // register wci_reqERR_5
  reg [2 : 0] wci_reqERR_5;
  wire [2 : 0] wci_reqERR_5$D_IN;
  wire wci_reqERR_5$EN;

  // register wci_reqERR_6
  reg [2 : 0] wci_reqERR_6;
  wire [2 : 0] wci_reqERR_6$D_IN;
  wire wci_reqERR_6$EN;

  // register wci_reqERR_7
  reg [2 : 0] wci_reqERR_7;
  wire [2 : 0] wci_reqERR_7$D_IN;
  wire wci_reqERR_7$EN;

  // register wci_reqERR_8
  reg [2 : 0] wci_reqERR_8;
  wire [2 : 0] wci_reqERR_8$D_IN;
  wire wci_reqERR_8$EN;

  // register wci_reqERR_9
  reg [2 : 0] wci_reqERR_9;
  wire [2 : 0] wci_reqERR_9$D_IN;
  wire wci_reqERR_9$EN;

  // register wci_reqFAIL
  reg [2 : 0] wci_reqFAIL;
  wire [2 : 0] wci_reqFAIL$D_IN;
  wire wci_reqFAIL$EN;

  // register wci_reqFAIL_1
  reg [2 : 0] wci_reqFAIL_1;
  wire [2 : 0] wci_reqFAIL_1$D_IN;
  wire wci_reqFAIL_1$EN;

  // register wci_reqFAIL_10
  reg [2 : 0] wci_reqFAIL_10;
  wire [2 : 0] wci_reqFAIL_10$D_IN;
  wire wci_reqFAIL_10$EN;

  // register wci_reqFAIL_11
  reg [2 : 0] wci_reqFAIL_11;
  wire [2 : 0] wci_reqFAIL_11$D_IN;
  wire wci_reqFAIL_11$EN;

  // register wci_reqFAIL_12
  reg [2 : 0] wci_reqFAIL_12;
  wire [2 : 0] wci_reqFAIL_12$D_IN;
  wire wci_reqFAIL_12$EN;

  // register wci_reqFAIL_13
  reg [2 : 0] wci_reqFAIL_13;
  wire [2 : 0] wci_reqFAIL_13$D_IN;
  wire wci_reqFAIL_13$EN;

  // register wci_reqFAIL_14
  reg [2 : 0] wci_reqFAIL_14;
  wire [2 : 0] wci_reqFAIL_14$D_IN;
  wire wci_reqFAIL_14$EN;

  // register wci_reqFAIL_2
  reg [2 : 0] wci_reqFAIL_2;
  wire [2 : 0] wci_reqFAIL_2$D_IN;
  wire wci_reqFAIL_2$EN;

  // register wci_reqFAIL_3
  reg [2 : 0] wci_reqFAIL_3;
  wire [2 : 0] wci_reqFAIL_3$D_IN;
  wire wci_reqFAIL_3$EN;

  // register wci_reqFAIL_4
  reg [2 : 0] wci_reqFAIL_4;
  wire [2 : 0] wci_reqFAIL_4$D_IN;
  wire wci_reqFAIL_4$EN;

  // register wci_reqFAIL_5
  reg [2 : 0] wci_reqFAIL_5;
  wire [2 : 0] wci_reqFAIL_5$D_IN;
  wire wci_reqFAIL_5$EN;

  // register wci_reqFAIL_6
  reg [2 : 0] wci_reqFAIL_6;
  wire [2 : 0] wci_reqFAIL_6$D_IN;
  wire wci_reqFAIL_6$EN;

  // register wci_reqFAIL_7
  reg [2 : 0] wci_reqFAIL_7;
  wire [2 : 0] wci_reqFAIL_7$D_IN;
  wire wci_reqFAIL_7$EN;

  // register wci_reqFAIL_8
  reg [2 : 0] wci_reqFAIL_8;
  wire [2 : 0] wci_reqFAIL_8$D_IN;
  wire wci_reqFAIL_8$EN;

  // register wci_reqFAIL_9
  reg [2 : 0] wci_reqFAIL_9;
  wire [2 : 0] wci_reqFAIL_9$D_IN;
  wire wci_reqFAIL_9$EN;

  // register wci_reqF_10_c_r
  reg wci_reqF_10_c_r;
  wire wci_reqF_10_c_r$D_IN, wci_reqF_10_c_r$EN;

  // register wci_reqF_10_q_0
  reg [71 : 0] wci_reqF_10_q_0;
  reg [71 : 0] wci_reqF_10_q_0$D_IN;
  wire wci_reqF_10_q_0$EN;

  // register wci_reqF_11_c_r
  reg wci_reqF_11_c_r;
  wire wci_reqF_11_c_r$D_IN, wci_reqF_11_c_r$EN;

  // register wci_reqF_11_q_0
  reg [71 : 0] wci_reqF_11_q_0;
  reg [71 : 0] wci_reqF_11_q_0$D_IN;
  wire wci_reqF_11_q_0$EN;

  // register wci_reqF_12_c_r
  reg wci_reqF_12_c_r;
  wire wci_reqF_12_c_r$D_IN, wci_reqF_12_c_r$EN;

  // register wci_reqF_12_q_0
  reg [71 : 0] wci_reqF_12_q_0;
  reg [71 : 0] wci_reqF_12_q_0$D_IN;
  wire wci_reqF_12_q_0$EN;

  // register wci_reqF_13_c_r
  reg wci_reqF_13_c_r;
  wire wci_reqF_13_c_r$D_IN, wci_reqF_13_c_r$EN;

  // register wci_reqF_13_q_0
  reg [71 : 0] wci_reqF_13_q_0;
  reg [71 : 0] wci_reqF_13_q_0$D_IN;
  wire wci_reqF_13_q_0$EN;

  // register wci_reqF_14_c_r
  reg wci_reqF_14_c_r;
  wire wci_reqF_14_c_r$D_IN, wci_reqF_14_c_r$EN;

  // register wci_reqF_14_q_0
  reg [71 : 0] wci_reqF_14_q_0;
  reg [71 : 0] wci_reqF_14_q_0$D_IN;
  wire wci_reqF_14_q_0$EN;

  // register wci_reqF_1_c_r
  reg wci_reqF_1_c_r;
  wire wci_reqF_1_c_r$D_IN, wci_reqF_1_c_r$EN;

  // register wci_reqF_1_q_0
  reg [71 : 0] wci_reqF_1_q_0;
  reg [71 : 0] wci_reqF_1_q_0$D_IN;
  wire wci_reqF_1_q_0$EN;

  // register wci_reqF_2_c_r
  reg wci_reqF_2_c_r;
  wire wci_reqF_2_c_r$D_IN, wci_reqF_2_c_r$EN;

  // register wci_reqF_2_q_0
  reg [71 : 0] wci_reqF_2_q_0;
  reg [71 : 0] wci_reqF_2_q_0$D_IN;
  wire wci_reqF_2_q_0$EN;

  // register wci_reqF_3_c_r
  reg wci_reqF_3_c_r;
  wire wci_reqF_3_c_r$D_IN, wci_reqF_3_c_r$EN;

  // register wci_reqF_3_q_0
  reg [71 : 0] wci_reqF_3_q_0;
  reg [71 : 0] wci_reqF_3_q_0$D_IN;
  wire wci_reqF_3_q_0$EN;

  // register wci_reqF_4_c_r
  reg wci_reqF_4_c_r;
  wire wci_reqF_4_c_r$D_IN, wci_reqF_4_c_r$EN;

  // register wci_reqF_4_q_0
  reg [71 : 0] wci_reqF_4_q_0;
  reg [71 : 0] wci_reqF_4_q_0$D_IN;
  wire wci_reqF_4_q_0$EN;

  // register wci_reqF_5_c_r
  reg wci_reqF_5_c_r;
  wire wci_reqF_5_c_r$D_IN, wci_reqF_5_c_r$EN;

  // register wci_reqF_5_q_0
  reg [71 : 0] wci_reqF_5_q_0;
  reg [71 : 0] wci_reqF_5_q_0$D_IN;
  wire wci_reqF_5_q_0$EN;

  // register wci_reqF_6_c_r
  reg wci_reqF_6_c_r;
  wire wci_reqF_6_c_r$D_IN, wci_reqF_6_c_r$EN;

  // register wci_reqF_6_q_0
  reg [71 : 0] wci_reqF_6_q_0;
  reg [71 : 0] wci_reqF_6_q_0$D_IN;
  wire wci_reqF_6_q_0$EN;

  // register wci_reqF_7_c_r
  reg wci_reqF_7_c_r;
  wire wci_reqF_7_c_r$D_IN, wci_reqF_7_c_r$EN;

  // register wci_reqF_7_q_0
  reg [71 : 0] wci_reqF_7_q_0;
  reg [71 : 0] wci_reqF_7_q_0$D_IN;
  wire wci_reqF_7_q_0$EN;

  // register wci_reqF_8_c_r
  reg wci_reqF_8_c_r;
  wire wci_reqF_8_c_r$D_IN, wci_reqF_8_c_r$EN;

  // register wci_reqF_8_q_0
  reg [71 : 0] wci_reqF_8_q_0;
  reg [71 : 0] wci_reqF_8_q_0$D_IN;
  wire wci_reqF_8_q_0$EN;

  // register wci_reqF_9_c_r
  reg wci_reqF_9_c_r;
  wire wci_reqF_9_c_r$D_IN, wci_reqF_9_c_r$EN;

  // register wci_reqF_9_q_0
  reg [71 : 0] wci_reqF_9_q_0;
  reg [71 : 0] wci_reqF_9_q_0$D_IN;
  wire wci_reqF_9_q_0$EN;

  // register wci_reqF_c_r
  reg wci_reqF_c_r;
  wire wci_reqF_c_r$D_IN, wci_reqF_c_r$EN;

  // register wci_reqF_q_0
  reg [71 : 0] wci_reqF_q_0;
  reg [71 : 0] wci_reqF_q_0$D_IN;
  wire wci_reqF_q_0$EN;

  // register wci_reqPend
  reg [1 : 0] wci_reqPend;
  reg [1 : 0] wci_reqPend$D_IN;
  wire wci_reqPend$EN;

  // register wci_reqPend_1
  reg [1 : 0] wci_reqPend_1;
  reg [1 : 0] wci_reqPend_1$D_IN;
  wire wci_reqPend_1$EN;

  // register wci_reqPend_10
  reg [1 : 0] wci_reqPend_10;
  reg [1 : 0] wci_reqPend_10$D_IN;
  wire wci_reqPend_10$EN;

  // register wci_reqPend_11
  reg [1 : 0] wci_reqPend_11;
  reg [1 : 0] wci_reqPend_11$D_IN;
  wire wci_reqPend_11$EN;

  // register wci_reqPend_12
  reg [1 : 0] wci_reqPend_12;
  reg [1 : 0] wci_reqPend_12$D_IN;
  wire wci_reqPend_12$EN;

  // register wci_reqPend_13
  reg [1 : 0] wci_reqPend_13;
  reg [1 : 0] wci_reqPend_13$D_IN;
  wire wci_reqPend_13$EN;

  // register wci_reqPend_14
  reg [1 : 0] wci_reqPend_14;
  reg [1 : 0] wci_reqPend_14$D_IN;
  wire wci_reqPend_14$EN;

  // register wci_reqPend_2
  reg [1 : 0] wci_reqPend_2;
  reg [1 : 0] wci_reqPend_2$D_IN;
  wire wci_reqPend_2$EN;

  // register wci_reqPend_3
  reg [1 : 0] wci_reqPend_3;
  reg [1 : 0] wci_reqPend_3$D_IN;
  wire wci_reqPend_3$EN;

  // register wci_reqPend_4
  reg [1 : 0] wci_reqPend_4;
  reg [1 : 0] wci_reqPend_4$D_IN;
  wire wci_reqPend_4$EN;

  // register wci_reqPend_5
  reg [1 : 0] wci_reqPend_5;
  reg [1 : 0] wci_reqPend_5$D_IN;
  wire wci_reqPend_5$EN;

  // register wci_reqPend_6
  reg [1 : 0] wci_reqPend_6;
  reg [1 : 0] wci_reqPend_6$D_IN;
  wire wci_reqPend_6$EN;

  // register wci_reqPend_7
  reg [1 : 0] wci_reqPend_7;
  reg [1 : 0] wci_reqPend_7$D_IN;
  wire wci_reqPend_7$EN;

  // register wci_reqPend_8
  reg [1 : 0] wci_reqPend_8;
  reg [1 : 0] wci_reqPend_8$D_IN;
  wire wci_reqPend_8$EN;

  // register wci_reqPend_9
  reg [1 : 0] wci_reqPend_9;
  reg [1 : 0] wci_reqPend_9$D_IN;
  wire wci_reqPend_9$EN;

  // register wci_reqTO
  reg [2 : 0] wci_reqTO;
  wire [2 : 0] wci_reqTO$D_IN;
  wire wci_reqTO$EN;

  // register wci_reqTO_1
  reg [2 : 0] wci_reqTO_1;
  wire [2 : 0] wci_reqTO_1$D_IN;
  wire wci_reqTO_1$EN;

  // register wci_reqTO_10
  reg [2 : 0] wci_reqTO_10;
  wire [2 : 0] wci_reqTO_10$D_IN;
  wire wci_reqTO_10$EN;

  // register wci_reqTO_11
  reg [2 : 0] wci_reqTO_11;
  wire [2 : 0] wci_reqTO_11$D_IN;
  wire wci_reqTO_11$EN;

  // register wci_reqTO_12
  reg [2 : 0] wci_reqTO_12;
  wire [2 : 0] wci_reqTO_12$D_IN;
  wire wci_reqTO_12$EN;

  // register wci_reqTO_13
  reg [2 : 0] wci_reqTO_13;
  wire [2 : 0] wci_reqTO_13$D_IN;
  wire wci_reqTO_13$EN;

  // register wci_reqTO_14
  reg [2 : 0] wci_reqTO_14;
  wire [2 : 0] wci_reqTO_14$D_IN;
  wire wci_reqTO_14$EN;

  // register wci_reqTO_2
  reg [2 : 0] wci_reqTO_2;
  wire [2 : 0] wci_reqTO_2$D_IN;
  wire wci_reqTO_2$EN;

  // register wci_reqTO_3
  reg [2 : 0] wci_reqTO_3;
  wire [2 : 0] wci_reqTO_3$D_IN;
  wire wci_reqTO_3$EN;

  // register wci_reqTO_4
  reg [2 : 0] wci_reqTO_4;
  wire [2 : 0] wci_reqTO_4$D_IN;
  wire wci_reqTO_4$EN;

  // register wci_reqTO_5
  reg [2 : 0] wci_reqTO_5;
  wire [2 : 0] wci_reqTO_5$D_IN;
  wire wci_reqTO_5$EN;

  // register wci_reqTO_6
  reg [2 : 0] wci_reqTO_6;
  wire [2 : 0] wci_reqTO_6$D_IN;
  wire wci_reqTO_6$EN;

  // register wci_reqTO_7
  reg [2 : 0] wci_reqTO_7;
  wire [2 : 0] wci_reqTO_7$D_IN;
  wire wci_reqTO_7$EN;

  // register wci_reqTO_8
  reg [2 : 0] wci_reqTO_8;
  wire [2 : 0] wci_reqTO_8$D_IN;
  wire wci_reqTO_8$EN;

  // register wci_reqTO_9
  reg [2 : 0] wci_reqTO_9;
  wire [2 : 0] wci_reqTO_9$D_IN;
  wire wci_reqTO_9$EN;

  // register wci_respTimr
  reg [31 : 0] wci_respTimr;
  wire [31 : 0] wci_respTimr$D_IN;
  wire wci_respTimr$EN;

  // register wci_respTimrAct
  reg wci_respTimrAct;
  wire wci_respTimrAct$D_IN, wci_respTimrAct$EN;

  // register wci_respTimrAct_1
  reg wci_respTimrAct_1;
  wire wci_respTimrAct_1$D_IN, wci_respTimrAct_1$EN;

  // register wci_respTimrAct_10
  reg wci_respTimrAct_10;
  wire wci_respTimrAct_10$D_IN, wci_respTimrAct_10$EN;

  // register wci_respTimrAct_11
  reg wci_respTimrAct_11;
  wire wci_respTimrAct_11$D_IN, wci_respTimrAct_11$EN;

  // register wci_respTimrAct_12
  reg wci_respTimrAct_12;
  wire wci_respTimrAct_12$D_IN, wci_respTimrAct_12$EN;

  // register wci_respTimrAct_13
  reg wci_respTimrAct_13;
  wire wci_respTimrAct_13$D_IN, wci_respTimrAct_13$EN;

  // register wci_respTimrAct_14
  reg wci_respTimrAct_14;
  wire wci_respTimrAct_14$D_IN, wci_respTimrAct_14$EN;

  // register wci_respTimrAct_2
  reg wci_respTimrAct_2;
  wire wci_respTimrAct_2$D_IN, wci_respTimrAct_2$EN;

  // register wci_respTimrAct_3
  reg wci_respTimrAct_3;
  wire wci_respTimrAct_3$D_IN, wci_respTimrAct_3$EN;

  // register wci_respTimrAct_4
  reg wci_respTimrAct_4;
  wire wci_respTimrAct_4$D_IN, wci_respTimrAct_4$EN;

  // register wci_respTimrAct_5
  reg wci_respTimrAct_5;
  wire wci_respTimrAct_5$D_IN, wci_respTimrAct_5$EN;

  // register wci_respTimrAct_6
  reg wci_respTimrAct_6;
  wire wci_respTimrAct_6$D_IN, wci_respTimrAct_6$EN;

  // register wci_respTimrAct_7
  reg wci_respTimrAct_7;
  wire wci_respTimrAct_7$D_IN, wci_respTimrAct_7$EN;

  // register wci_respTimrAct_8
  reg wci_respTimrAct_8;
  wire wci_respTimrAct_8$D_IN, wci_respTimrAct_8$EN;

  // register wci_respTimrAct_9
  reg wci_respTimrAct_9;
  wire wci_respTimrAct_9$D_IN, wci_respTimrAct_9$EN;

  // register wci_respTimr_1
  reg [31 : 0] wci_respTimr_1;
  wire [31 : 0] wci_respTimr_1$D_IN;
  wire wci_respTimr_1$EN;

  // register wci_respTimr_10
  reg [31 : 0] wci_respTimr_10;
  wire [31 : 0] wci_respTimr_10$D_IN;
  wire wci_respTimr_10$EN;

  // register wci_respTimr_11
  reg [31 : 0] wci_respTimr_11;
  wire [31 : 0] wci_respTimr_11$D_IN;
  wire wci_respTimr_11$EN;

  // register wci_respTimr_12
  reg [31 : 0] wci_respTimr_12;
  wire [31 : 0] wci_respTimr_12$D_IN;
  wire wci_respTimr_12$EN;

  // register wci_respTimr_13
  reg [31 : 0] wci_respTimr_13;
  wire [31 : 0] wci_respTimr_13$D_IN;
  wire wci_respTimr_13$EN;

  // register wci_respTimr_14
  reg [31 : 0] wci_respTimr_14;
  wire [31 : 0] wci_respTimr_14$D_IN;
  wire wci_respTimr_14$EN;

  // register wci_respTimr_2
  reg [31 : 0] wci_respTimr_2;
  wire [31 : 0] wci_respTimr_2$D_IN;
  wire wci_respTimr_2$EN;

  // register wci_respTimr_3
  reg [31 : 0] wci_respTimr_3;
  wire [31 : 0] wci_respTimr_3$D_IN;
  wire wci_respTimr_3$EN;

  // register wci_respTimr_4
  reg [31 : 0] wci_respTimr_4;
  wire [31 : 0] wci_respTimr_4$D_IN;
  wire wci_respTimr_4$EN;

  // register wci_respTimr_5
  reg [31 : 0] wci_respTimr_5;
  wire [31 : 0] wci_respTimr_5$D_IN;
  wire wci_respTimr_5$EN;

  // register wci_respTimr_6
  reg [31 : 0] wci_respTimr_6;
  wire [31 : 0] wci_respTimr_6$D_IN;
  wire wci_respTimr_6$EN;

  // register wci_respTimr_7
  reg [31 : 0] wci_respTimr_7;
  wire [31 : 0] wci_respTimr_7$D_IN;
  wire wci_respTimr_7$EN;

  // register wci_respTimr_8
  reg [31 : 0] wci_respTimr_8;
  wire [31 : 0] wci_respTimr_8$D_IN;
  wire wci_respTimr_8$EN;

  // register wci_respTimr_9
  reg [31 : 0] wci_respTimr_9;
  wire [31 : 0] wci_respTimr_9$D_IN;
  wire wci_respTimr_9$EN;

  // register wci_sThreadBusy_d
  reg wci_sThreadBusy_d;
  wire wci_sThreadBusy_d$D_IN, wci_sThreadBusy_d$EN;

  // register wci_sThreadBusy_d_1
  reg wci_sThreadBusy_d_1;
  wire wci_sThreadBusy_d_1$D_IN, wci_sThreadBusy_d_1$EN;

  // register wci_sThreadBusy_d_10
  reg wci_sThreadBusy_d_10;
  wire wci_sThreadBusy_d_10$D_IN, wci_sThreadBusy_d_10$EN;

  // register wci_sThreadBusy_d_11
  reg wci_sThreadBusy_d_11;
  wire wci_sThreadBusy_d_11$D_IN, wci_sThreadBusy_d_11$EN;

  // register wci_sThreadBusy_d_12
  reg wci_sThreadBusy_d_12;
  wire wci_sThreadBusy_d_12$D_IN, wci_sThreadBusy_d_12$EN;

  // register wci_sThreadBusy_d_13
  reg wci_sThreadBusy_d_13;
  wire wci_sThreadBusy_d_13$D_IN, wci_sThreadBusy_d_13$EN;

  // register wci_sThreadBusy_d_14
  reg wci_sThreadBusy_d_14;
  wire wci_sThreadBusy_d_14$D_IN, wci_sThreadBusy_d_14$EN;

  // register wci_sThreadBusy_d_2
  reg wci_sThreadBusy_d_2;
  wire wci_sThreadBusy_d_2$D_IN, wci_sThreadBusy_d_2$EN;

  // register wci_sThreadBusy_d_3
  reg wci_sThreadBusy_d_3;
  wire wci_sThreadBusy_d_3$D_IN, wci_sThreadBusy_d_3$EN;

  // register wci_sThreadBusy_d_4
  reg wci_sThreadBusy_d_4;
  wire wci_sThreadBusy_d_4$D_IN, wci_sThreadBusy_d_4$EN;

  // register wci_sThreadBusy_d_5
  reg wci_sThreadBusy_d_5;
  wire wci_sThreadBusy_d_5$D_IN, wci_sThreadBusy_d_5$EN;

  // register wci_sThreadBusy_d_6
  reg wci_sThreadBusy_d_6;
  wire wci_sThreadBusy_d_6$D_IN, wci_sThreadBusy_d_6$EN;

  // register wci_sThreadBusy_d_7
  reg wci_sThreadBusy_d_7;
  wire wci_sThreadBusy_d_7$D_IN, wci_sThreadBusy_d_7$EN;

  // register wci_sThreadBusy_d_8
  reg wci_sThreadBusy_d_8;
  wire wci_sThreadBusy_d_8$D_IN, wci_sThreadBusy_d_8$EN;

  // register wci_sThreadBusy_d_9
  reg wci_sThreadBusy_d_9;
  wire wci_sThreadBusy_d_9$D_IN, wci_sThreadBusy_d_9$EN;

  // register wci_sfCap
  reg wci_sfCap;
  wire wci_sfCap$D_IN, wci_sfCap$EN;

  // register wci_sfCapClear
  reg wci_sfCapClear;
  wire wci_sfCapClear$D_IN, wci_sfCapClear$EN;

  // register wci_sfCapClear_10
  reg wci_sfCapClear_10;
  wire wci_sfCapClear_10$D_IN, wci_sfCapClear_10$EN;

  // register wci_sfCapClear_11
  reg wci_sfCapClear_11;
  wire wci_sfCapClear_11$D_IN, wci_sfCapClear_11$EN;

  // register wci_sfCapClear_12
  reg wci_sfCapClear_12;
  wire wci_sfCapClear_12$D_IN, wci_sfCapClear_12$EN;

  // register wci_sfCapClear_13
  reg wci_sfCapClear_13;
  wire wci_sfCapClear_13$D_IN, wci_sfCapClear_13$EN;

  // register wci_sfCapClear_14
  reg wci_sfCapClear_14;
  wire wci_sfCapClear_14$D_IN, wci_sfCapClear_14$EN;

  // register wci_sfCapClear_1_1
  reg wci_sfCapClear_1_1;
  wire wci_sfCapClear_1_1$D_IN, wci_sfCapClear_1_1$EN;

  // register wci_sfCapClear_2
  reg wci_sfCapClear_2;
  wire wci_sfCapClear_2$D_IN, wci_sfCapClear_2$EN;

  // register wci_sfCapClear_3
  reg wci_sfCapClear_3;
  wire wci_sfCapClear_3$D_IN, wci_sfCapClear_3$EN;

  // register wci_sfCapClear_4
  reg wci_sfCapClear_4;
  wire wci_sfCapClear_4$D_IN, wci_sfCapClear_4$EN;

  // register wci_sfCapClear_5
  reg wci_sfCapClear_5;
  wire wci_sfCapClear_5$D_IN, wci_sfCapClear_5$EN;

  // register wci_sfCapClear_6
  reg wci_sfCapClear_6;
  wire wci_sfCapClear_6$D_IN, wci_sfCapClear_6$EN;

  // register wci_sfCapClear_7
  reg wci_sfCapClear_7;
  wire wci_sfCapClear_7$D_IN, wci_sfCapClear_7$EN;

  // register wci_sfCapClear_8
  reg wci_sfCapClear_8;
  wire wci_sfCapClear_8$D_IN, wci_sfCapClear_8$EN;

  // register wci_sfCapClear_9
  reg wci_sfCapClear_9;
  wire wci_sfCapClear_9$D_IN, wci_sfCapClear_9$EN;

  // register wci_sfCapSet
  reg wci_sfCapSet;
  wire wci_sfCapSet$D_IN, wci_sfCapSet$EN;

  // register wci_sfCapSet_10
  reg wci_sfCapSet_10;
  wire wci_sfCapSet_10$D_IN, wci_sfCapSet_10$EN;

  // register wci_sfCapSet_11
  reg wci_sfCapSet_11;
  wire wci_sfCapSet_11$D_IN, wci_sfCapSet_11$EN;

  // register wci_sfCapSet_12
  reg wci_sfCapSet_12;
  wire wci_sfCapSet_12$D_IN, wci_sfCapSet_12$EN;

  // register wci_sfCapSet_13
  reg wci_sfCapSet_13;
  wire wci_sfCapSet_13$D_IN, wci_sfCapSet_13$EN;

  // register wci_sfCapSet_14
  reg wci_sfCapSet_14;
  wire wci_sfCapSet_14$D_IN, wci_sfCapSet_14$EN;

  // register wci_sfCapSet_1_1
  reg wci_sfCapSet_1_1;
  wire wci_sfCapSet_1_1$D_IN, wci_sfCapSet_1_1$EN;

  // register wci_sfCapSet_2
  reg wci_sfCapSet_2;
  wire wci_sfCapSet_2$D_IN, wci_sfCapSet_2$EN;

  // register wci_sfCapSet_3
  reg wci_sfCapSet_3;
  wire wci_sfCapSet_3$D_IN, wci_sfCapSet_3$EN;

  // register wci_sfCapSet_4
  reg wci_sfCapSet_4;
  wire wci_sfCapSet_4$D_IN, wci_sfCapSet_4$EN;

  // register wci_sfCapSet_5
  reg wci_sfCapSet_5;
  wire wci_sfCapSet_5$D_IN, wci_sfCapSet_5$EN;

  // register wci_sfCapSet_6
  reg wci_sfCapSet_6;
  wire wci_sfCapSet_6$D_IN, wci_sfCapSet_6$EN;

  // register wci_sfCapSet_7
  reg wci_sfCapSet_7;
  wire wci_sfCapSet_7$D_IN, wci_sfCapSet_7$EN;

  // register wci_sfCapSet_8
  reg wci_sfCapSet_8;
  wire wci_sfCapSet_8$D_IN, wci_sfCapSet_8$EN;

  // register wci_sfCapSet_9
  reg wci_sfCapSet_9;
  wire wci_sfCapSet_9$D_IN, wci_sfCapSet_9$EN;

  // register wci_sfCap_1
  reg wci_sfCap_1;
  wire wci_sfCap_1$D_IN, wci_sfCap_1$EN;

  // register wci_sfCap_10
  reg wci_sfCap_10;
  wire wci_sfCap_10$D_IN, wci_sfCap_10$EN;

  // register wci_sfCap_11
  reg wci_sfCap_11;
  wire wci_sfCap_11$D_IN, wci_sfCap_11$EN;

  // register wci_sfCap_12
  reg wci_sfCap_12;
  wire wci_sfCap_12$D_IN, wci_sfCap_12$EN;

  // register wci_sfCap_13
  reg wci_sfCap_13;
  wire wci_sfCap_13$D_IN, wci_sfCap_13$EN;

  // register wci_sfCap_14
  reg wci_sfCap_14;
  wire wci_sfCap_14$D_IN, wci_sfCap_14$EN;

  // register wci_sfCap_2
  reg wci_sfCap_2;
  wire wci_sfCap_2$D_IN, wci_sfCap_2$EN;

  // register wci_sfCap_3
  reg wci_sfCap_3;
  wire wci_sfCap_3$D_IN, wci_sfCap_3$EN;

  // register wci_sfCap_4
  reg wci_sfCap_4;
  wire wci_sfCap_4$D_IN, wci_sfCap_4$EN;

  // register wci_sfCap_5
  reg wci_sfCap_5;
  wire wci_sfCap_5$D_IN, wci_sfCap_5$EN;

  // register wci_sfCap_6
  reg wci_sfCap_6;
  wire wci_sfCap_6$D_IN, wci_sfCap_6$EN;

  // register wci_sfCap_7
  reg wci_sfCap_7;
  wire wci_sfCap_7$D_IN, wci_sfCap_7$EN;

  // register wci_sfCap_8
  reg wci_sfCap_8;
  wire wci_sfCap_8$D_IN, wci_sfCap_8$EN;

  // register wci_sfCap_9
  reg wci_sfCap_9;
  wire wci_sfCap_9$D_IN, wci_sfCap_9$EN;

  // register wci_slvPresent
  reg wci_slvPresent;
  wire wci_slvPresent$D_IN, wci_slvPresent$EN;

  // register wci_slvPresent_1
  reg wci_slvPresent_1;
  wire wci_slvPresent_1$D_IN, wci_slvPresent_1$EN;

  // register wci_slvPresent_10
  reg wci_slvPresent_10;
  wire wci_slvPresent_10$D_IN, wci_slvPresent_10$EN;

  // register wci_slvPresent_11
  reg wci_slvPresent_11;
  wire wci_slvPresent_11$D_IN, wci_slvPresent_11$EN;

  // register wci_slvPresent_12
  reg wci_slvPresent_12;
  wire wci_slvPresent_12$D_IN, wci_slvPresent_12$EN;

  // register wci_slvPresent_13
  reg wci_slvPresent_13;
  wire wci_slvPresent_13$D_IN, wci_slvPresent_13$EN;

  // register wci_slvPresent_14
  reg wci_slvPresent_14;
  wire wci_slvPresent_14$D_IN, wci_slvPresent_14$EN;

  // register wci_slvPresent_2
  reg wci_slvPresent_2;
  wire wci_slvPresent_2$D_IN, wci_slvPresent_2$EN;

  // register wci_slvPresent_3
  reg wci_slvPresent_3;
  wire wci_slvPresent_3$D_IN, wci_slvPresent_3$EN;

  // register wci_slvPresent_4
  reg wci_slvPresent_4;
  wire wci_slvPresent_4$D_IN, wci_slvPresent_4$EN;

  // register wci_slvPresent_5
  reg wci_slvPresent_5;
  wire wci_slvPresent_5$D_IN, wci_slvPresent_5$EN;

  // register wci_slvPresent_6
  reg wci_slvPresent_6;
  wire wci_slvPresent_6$D_IN, wci_slvPresent_6$EN;

  // register wci_slvPresent_7
  reg wci_slvPresent_7;
  wire wci_slvPresent_7$D_IN, wci_slvPresent_7$EN;

  // register wci_slvPresent_8
  reg wci_slvPresent_8;
  wire wci_slvPresent_8$D_IN, wci_slvPresent_8$EN;

  // register wci_slvPresent_9
  reg wci_slvPresent_9;
  wire wci_slvPresent_9$D_IN, wci_slvPresent_9$EN;

  // register wci_wReset_n
  reg wci_wReset_n;
  wire wci_wReset_n$D_IN, wci_wReset_n$EN;

  // register wci_wReset_n_1
  reg wci_wReset_n_1;
  wire wci_wReset_n_1$D_IN, wci_wReset_n_1$EN;

  // register wci_wReset_n_10
  reg wci_wReset_n_10;
  wire wci_wReset_n_10$D_IN, wci_wReset_n_10$EN;

  // register wci_wReset_n_11
  reg wci_wReset_n_11;
  wire wci_wReset_n_11$D_IN, wci_wReset_n_11$EN;

  // register wci_wReset_n_12
  reg wci_wReset_n_12;
  wire wci_wReset_n_12$D_IN, wci_wReset_n_12$EN;

  // register wci_wReset_n_13
  reg wci_wReset_n_13;
  wire wci_wReset_n_13$D_IN, wci_wReset_n_13$EN;

  // register wci_wReset_n_14
  reg wci_wReset_n_14;
  wire wci_wReset_n_14$D_IN, wci_wReset_n_14$EN;

  // register wci_wReset_n_2
  reg wci_wReset_n_2;
  wire wci_wReset_n_2$D_IN, wci_wReset_n_2$EN;

  // register wci_wReset_n_3
  reg wci_wReset_n_3;
  wire wci_wReset_n_3$D_IN, wci_wReset_n_3$EN;

  // register wci_wReset_n_4
  reg wci_wReset_n_4;
  wire wci_wReset_n_4$D_IN, wci_wReset_n_4$EN;

  // register wci_wReset_n_5
  reg wci_wReset_n_5;
  wire wci_wReset_n_5$D_IN, wci_wReset_n_5$EN;

  // register wci_wReset_n_6
  reg wci_wReset_n_6;
  wire wci_wReset_n_6$D_IN, wci_wReset_n_6$EN;

  // register wci_wReset_n_7
  reg wci_wReset_n_7;
  wire wci_wReset_n_7$D_IN, wci_wReset_n_7$EN;

  // register wci_wReset_n_8
  reg wci_wReset_n_8;
  wire wci_wReset_n_8$D_IN, wci_wReset_n_8$EN;

  // register wci_wReset_n_9
  reg wci_wReset_n_9;
  wire wci_wReset_n_9$D_IN, wci_wReset_n_9$EN;

  // register wci_wStatus
  reg [31 : 0] wci_wStatus;
  wire [31 : 0] wci_wStatus$D_IN;
  wire wci_wStatus$EN;

  // register wci_wStatus_1
  reg [31 : 0] wci_wStatus_1;
  wire [31 : 0] wci_wStatus_1$D_IN;
  wire wci_wStatus_1$EN;

  // register wci_wStatus_10
  reg [31 : 0] wci_wStatus_10;
  wire [31 : 0] wci_wStatus_10$D_IN;
  wire wci_wStatus_10$EN;

  // register wci_wStatus_11
  reg [31 : 0] wci_wStatus_11;
  wire [31 : 0] wci_wStatus_11$D_IN;
  wire wci_wStatus_11$EN;

  // register wci_wStatus_12
  reg [31 : 0] wci_wStatus_12;
  wire [31 : 0] wci_wStatus_12$D_IN;
  wire wci_wStatus_12$EN;

  // register wci_wStatus_13
  reg [31 : 0] wci_wStatus_13;
  wire [31 : 0] wci_wStatus_13$D_IN;
  wire wci_wStatus_13$EN;

  // register wci_wStatus_14
  reg [31 : 0] wci_wStatus_14;
  wire [31 : 0] wci_wStatus_14$D_IN;
  wire wci_wStatus_14$EN;

  // register wci_wStatus_2
  reg [31 : 0] wci_wStatus_2;
  wire [31 : 0] wci_wStatus_2$D_IN;
  wire wci_wStatus_2$EN;

  // register wci_wStatus_3
  reg [31 : 0] wci_wStatus_3;
  wire [31 : 0] wci_wStatus_3$D_IN;
  wire wci_wStatus_3$EN;

  // register wci_wStatus_4
  reg [31 : 0] wci_wStatus_4;
  wire [31 : 0] wci_wStatus_4$D_IN;
  wire wci_wStatus_4$EN;

  // register wci_wStatus_5
  reg [31 : 0] wci_wStatus_5;
  wire [31 : 0] wci_wStatus_5$D_IN;
  wire wci_wStatus_5$EN;

  // register wci_wStatus_6
  reg [31 : 0] wci_wStatus_6;
  wire [31 : 0] wci_wStatus_6$D_IN;
  wire wci_wStatus_6$EN;

  // register wci_wStatus_7
  reg [31 : 0] wci_wStatus_7;
  wire [31 : 0] wci_wStatus_7$D_IN;
  wire wci_wStatus_7$EN;

  // register wci_wStatus_8
  reg [31 : 0] wci_wStatus_8;
  wire [31 : 0] wci_wStatus_8$D_IN;
  wire wci_wStatus_8$EN;

  // register wci_wStatus_9
  reg [31 : 0] wci_wStatus_9;
  wire [31 : 0] wci_wStatus_9$D_IN;
  wire wci_wStatus_9$EN;

  // register wci_wTimeout
  reg [4 : 0] wci_wTimeout;
  wire [4 : 0] wci_wTimeout$D_IN;
  wire wci_wTimeout$EN;

  // register wci_wTimeout_1
  reg [4 : 0] wci_wTimeout_1;
  wire [4 : 0] wci_wTimeout_1$D_IN;
  wire wci_wTimeout_1$EN;

  // register wci_wTimeout_10
  reg [4 : 0] wci_wTimeout_10;
  wire [4 : 0] wci_wTimeout_10$D_IN;
  wire wci_wTimeout_10$EN;

  // register wci_wTimeout_11
  reg [4 : 0] wci_wTimeout_11;
  wire [4 : 0] wci_wTimeout_11$D_IN;
  wire wci_wTimeout_11$EN;

  // register wci_wTimeout_12
  reg [4 : 0] wci_wTimeout_12;
  wire [4 : 0] wci_wTimeout_12$D_IN;
  wire wci_wTimeout_12$EN;

  // register wci_wTimeout_13
  reg [4 : 0] wci_wTimeout_13;
  wire [4 : 0] wci_wTimeout_13$D_IN;
  wire wci_wTimeout_13$EN;

  // register wci_wTimeout_14
  reg [4 : 0] wci_wTimeout_14;
  wire [4 : 0] wci_wTimeout_14$D_IN;
  wire wci_wTimeout_14$EN;

  // register wci_wTimeout_2
  reg [4 : 0] wci_wTimeout_2;
  wire [4 : 0] wci_wTimeout_2$D_IN;
  wire wci_wTimeout_2$EN;

  // register wci_wTimeout_3
  reg [4 : 0] wci_wTimeout_3;
  wire [4 : 0] wci_wTimeout_3$D_IN;
  wire wci_wTimeout_3$EN;

  // register wci_wTimeout_4
  reg [4 : 0] wci_wTimeout_4;
  wire [4 : 0] wci_wTimeout_4$D_IN;
  wire wci_wTimeout_4$EN;

  // register wci_wTimeout_5
  reg [4 : 0] wci_wTimeout_5;
  wire [4 : 0] wci_wTimeout_5$D_IN;
  wire wci_wTimeout_5$EN;

  // register wci_wTimeout_6
  reg [4 : 0] wci_wTimeout_6;
  wire [4 : 0] wci_wTimeout_6$D_IN;
  wire wci_wTimeout_6$EN;

  // register wci_wTimeout_7
  reg [4 : 0] wci_wTimeout_7;
  wire [4 : 0] wci_wTimeout_7$D_IN;
  wire wci_wTimeout_7$EN;

  // register wci_wTimeout_8
  reg [4 : 0] wci_wTimeout_8;
  wire [4 : 0] wci_wTimeout_8$D_IN;
  wire wci_wTimeout_8$EN;

  // register wci_wTimeout_9
  reg [4 : 0] wci_wTimeout_9;
  wire [4 : 0] wci_wTimeout_9$D_IN;
  wire wci_wTimeout_9$EN;

  // register wrkAct
  reg [3 : 0] wrkAct;
  reg [3 : 0] wrkAct$D_IN;
  wire wrkAct$EN;

  // ports of submodule adminResp1F
  wire [32 : 0] adminResp1F$D_IN, adminResp1F$D_OUT;
  wire adminResp1F$CLR,
       adminResp1F$DEQ,
       adminResp1F$EMPTY_N,
       adminResp1F$ENQ,
       adminResp1F$FULL_N;

  // ports of submodule adminResp2F
  reg [32 : 0] adminResp2F$D_IN;
  wire [32 : 0] adminResp2F$D_OUT;
  wire adminResp2F$CLR,
       adminResp2F$DEQ,
       adminResp2F$EMPTY_N,
       adminResp2F$ENQ,
       adminResp2F$FULL_N;

  // ports of submodule adminResp3F
  wire [32 : 0] adminResp3F$D_IN, adminResp3F$D_OUT;
  wire adminResp3F$CLR,
       adminResp3F$DEQ,
       adminResp3F$EMPTY_N,
       adminResp3F$ENQ,
       adminResp3F$FULL_N;

  // ports of submodule adminResp4F
  wire [32 : 0] adminResp4F$D_IN, adminResp4F$D_OUT;
  wire adminResp4F$CLR,
       adminResp4F$DEQ,
       adminResp4F$EMPTY_N,
       adminResp4F$ENQ,
       adminResp4F$FULL_N;

  // ports of submodule adminRespF
  wire [32 : 0] adminRespF$D_IN, adminRespF$D_OUT;
  wire adminRespF$CLR,
       adminRespF$DEQ,
       adminRespF$EMPTY_N,
       adminRespF$ENQ,
       adminRespF$FULL_N;

  // ports of submodule cpReqF
  wire [58 : 0] cpReqF$D_IN, cpReqF$D_OUT;
  wire cpReqF$CLR, cpReqF$DEQ, cpReqF$EMPTY_N, cpReqF$ENQ, cpReqF$FULL_N;

  // ports of submodule cpRespF
  wire [39 : 0] cpRespF$D_IN, cpRespF$D_OUT;
  wire cpRespF$CLR, cpRespF$DEQ, cpRespF$EMPTY_N, cpRespF$ENQ, cpRespF$FULL_N;

`ifdef not
  // ports of submodule dna_dna
  wire dna_dna$CLK, dna_dna$DIN, dna_dna$DOUT, dna_dna$READ, dna_dna$SHIFT;

  // ports of submodule rom_memory
  wire [31 : 0] rom_memory$DI, rom_memory$DO;
  wire [9 : 0] rom_memory$ADDR;
  wire rom_memory$EN, rom_memory$WE;

  // ports of submodule rom_serverAdapter_outDataCore
  wire [31 : 0] rom_serverAdapter_outDataCore$D_IN,
		rom_serverAdapter_outDataCore$D_OUT;
  wire rom_serverAdapter_outDataCore$CLR,
       rom_serverAdapter_outDataCore$DEQ,
       rom_serverAdapter_outDataCore$EMPTY_N,
       rom_serverAdapter_outDataCore$ENQ,
       rom_serverAdapter_outDataCore$FULL_N;

  // ports of submodule timeServ_disableServo
  wire timeServ_disableServo$dD_OUT,
       timeServ_disableServo$sD_IN,
       timeServ_disableServo$sEN,
       timeServ_disableServo$sRDY;

  // ports of submodule timeServ_nowInCC
  wire [63 : 0] timeServ_nowInCC$dD_OUT, timeServ_nowInCC$sD_IN;
  wire timeServ_nowInCC$sEN, timeServ_nowInCC$sRDY;

  // ports of submodule timeServ_ppsDisablePPS
  wire timeServ_ppsDisablePPS$dD_OUT,
       timeServ_ppsDisablePPS$sD_IN,
       timeServ_ppsDisablePPS$sEN,
       timeServ_ppsDisablePPS$sRDY;

  // ports of submodule timeServ_ppsLostCC
  wire timeServ_ppsLostCC$dD_OUT,
       timeServ_ppsLostCC$sD_IN,
       timeServ_ppsLostCC$sEN,
       timeServ_ppsLostCC$sRDY;

  // ports of submodule timeServ_ppsOKCC
  wire timeServ_ppsOKCC$dD_OUT,
       timeServ_ppsOKCC$sD_IN,
       timeServ_ppsOKCC$sEN,
       timeServ_ppsOKCC$sRDY;

  // ports of submodule timeServ_ppsOutMode
  wire [1 : 0] timeServ_ppsOutMode$dD_OUT, timeServ_ppsOutMode$sD_IN;
  wire timeServ_ppsOutMode$sEN, timeServ_ppsOutMode$sRDY;

  // ports of submodule timeServ_refPerPPS
  wire [27 : 0] timeServ_refPerPPS$dD_OUT, timeServ_refPerPPS$sD_IN;
  wire timeServ_refPerPPS$sEN, timeServ_refPerPPS$sRDY;

  // ports of submodule timeServ_rollingPPSIn
  wire [7 : 0] timeServ_rollingPPSIn$dD_OUT, timeServ_rollingPPSIn$sD_IN;
  wire timeServ_rollingPPSIn$sEN, timeServ_rollingPPSIn$sRDY;

  // ports of submodule timeServ_setRefF
  wire [63 : 0] timeServ_setRefF$dD_OUT, timeServ_setRefF$sD_IN;
  wire timeServ_setRefF$dDEQ,
       timeServ_setRefF$dEMPTY_N,
       timeServ_setRefF$sENQ,
       timeServ_setRefF$sFULL_N;
`endif

  // ports of submodule wci_mReset
  wire wci_mReset$ASSERT_IN, wci_mReset$OUT_RST;

  // ports of submodule wci_mReset_1
  wire wci_mReset_1$ASSERT_IN, wci_mReset_1$OUT_RST;

  // ports of submodule wci_mReset_10
  wire wci_mReset_10$ASSERT_IN, wci_mReset_10$OUT_RST;

  // ports of submodule wci_mReset_11
  wire wci_mReset_11$ASSERT_IN, wci_mReset_11$OUT_RST;

  // ports of submodule wci_mReset_12
  wire wci_mReset_12$ASSERT_IN, wci_mReset_12$OUT_RST;

  // ports of submodule wci_mReset_13
  wire wci_mReset_13$ASSERT_IN, wci_mReset_13$OUT_RST;

  // ports of submodule wci_mReset_14
  wire wci_mReset_14$ASSERT_IN, wci_mReset_14$OUT_RST;

  // ports of submodule wci_mReset_2
  wire wci_mReset_2$ASSERT_IN, wci_mReset_2$OUT_RST;

  // ports of submodule wci_mReset_3
  wire wci_mReset_3$ASSERT_IN, wci_mReset_3$OUT_RST;

  // ports of submodule wci_mReset_4
  wire wci_mReset_4$ASSERT_IN, wci_mReset_4$OUT_RST;

  // ports of submodule wci_mReset_5
  wire wci_mReset_5$ASSERT_IN, wci_mReset_5$OUT_RST;

  // ports of submodule wci_mReset_6
  wire wci_mReset_6$ASSERT_IN, wci_mReset_6$OUT_RST;

  // ports of submodule wci_mReset_7
  wire wci_mReset_7$ASSERT_IN, wci_mReset_7$OUT_RST;

  // ports of submodule wci_mReset_8
  wire wci_mReset_8$ASSERT_IN, wci_mReset_8$OUT_RST;

  // ports of submodule wci_mReset_9
  wire wci_mReset_9$ASSERT_IN, wci_mReset_9$OUT_RST;

  // ports of submodule wci_respF
  reg [33 : 0] wci_respF$D_IN;
  wire [33 : 0] wci_respF$D_OUT;
  wire wci_respF$CLR,
       wci_respF$DEQ,
       wci_respF$EMPTY_N,
       wci_respF$ENQ,
       wci_respF$FULL_N;

  // ports of submodule wci_respF_1
  reg [33 : 0] wci_respF_1$D_IN;
  wire [33 : 0] wci_respF_1$D_OUT;
  wire wci_respF_1$CLR,
       wci_respF_1$DEQ,
       wci_respF_1$EMPTY_N,
       wci_respF_1$ENQ,
       wci_respF_1$FULL_N;

  // ports of submodule wci_respF_10
  reg [33 : 0] wci_respF_10$D_IN;
  wire [33 : 0] wci_respF_10$D_OUT;
  wire wci_respF_10$CLR,
       wci_respF_10$DEQ,
       wci_respF_10$EMPTY_N,
       wci_respF_10$ENQ,
       wci_respF_10$FULL_N;

  // ports of submodule wci_respF_11
  reg [33 : 0] wci_respF_11$D_IN;
  wire [33 : 0] wci_respF_11$D_OUT;
  wire wci_respF_11$CLR,
       wci_respF_11$DEQ,
       wci_respF_11$EMPTY_N,
       wci_respF_11$ENQ,
       wci_respF_11$FULL_N;

  // ports of submodule wci_respF_12
  reg [33 : 0] wci_respF_12$D_IN;
  wire [33 : 0] wci_respF_12$D_OUT;
  wire wci_respF_12$CLR,
       wci_respF_12$DEQ,
       wci_respF_12$EMPTY_N,
       wci_respF_12$ENQ,
       wci_respF_12$FULL_N;

  // ports of submodule wci_respF_13
  reg [33 : 0] wci_respF_13$D_IN;
  wire [33 : 0] wci_respF_13$D_OUT;
  wire wci_respF_13$CLR,
       wci_respF_13$DEQ,
       wci_respF_13$EMPTY_N,
       wci_respF_13$ENQ,
       wci_respF_13$FULL_N;

  // ports of submodule wci_respF_14
  reg [33 : 0] wci_respF_14$D_IN;
  wire [33 : 0] wci_respF_14$D_OUT;
  wire wci_respF_14$CLR,
       wci_respF_14$DEQ,
       wci_respF_14$EMPTY_N,
       wci_respF_14$ENQ,
       wci_respF_14$FULL_N;

  // ports of submodule wci_respF_2
  reg [33 : 0] wci_respF_2$D_IN;
  wire [33 : 0] wci_respF_2$D_OUT;
  wire wci_respF_2$CLR,
       wci_respF_2$DEQ,
       wci_respF_2$EMPTY_N,
       wci_respF_2$ENQ,
       wci_respF_2$FULL_N;

  // ports of submodule wci_respF_3
  reg [33 : 0] wci_respF_3$D_IN;
  wire [33 : 0] wci_respF_3$D_OUT;
  wire wci_respF_3$CLR,
       wci_respF_3$DEQ,
       wci_respF_3$EMPTY_N,
       wci_respF_3$ENQ,
       wci_respF_3$FULL_N;

  // ports of submodule wci_respF_4
  reg [33 : 0] wci_respF_4$D_IN;
  wire [33 : 0] wci_respF_4$D_OUT;
  wire wci_respF_4$CLR,
       wci_respF_4$DEQ,
       wci_respF_4$EMPTY_N,
       wci_respF_4$ENQ,
       wci_respF_4$FULL_N;

  // ports of submodule wci_respF_5
  reg [33 : 0] wci_respF_5$D_IN;
  wire [33 : 0] wci_respF_5$D_OUT;
  wire wci_respF_5$CLR,
       wci_respF_5$DEQ,
       wci_respF_5$EMPTY_N,
       wci_respF_5$ENQ,
       wci_respF_5$FULL_N;

  // ports of submodule wci_respF_6
  reg [33 : 0] wci_respF_6$D_IN;
  wire [33 : 0] wci_respF_6$D_OUT;
  wire wci_respF_6$CLR,
       wci_respF_6$DEQ,
       wci_respF_6$EMPTY_N,
       wci_respF_6$ENQ,
       wci_respF_6$FULL_N;

  // ports of submodule wci_respF_7
  reg [33 : 0] wci_respF_7$D_IN;
  wire [33 : 0] wci_respF_7$D_OUT;
  wire wci_respF_7$CLR,
       wci_respF_7$DEQ,
       wci_respF_7$EMPTY_N,
       wci_respF_7$ENQ,
       wci_respF_7$FULL_N;

  // ports of submodule wci_respF_8
  reg [33 : 0] wci_respF_8$D_IN;
  wire [33 : 0] wci_respF_8$D_OUT;
  wire wci_respF_8$CLR,
       wci_respF_8$DEQ,
       wci_respF_8$EMPTY_N,
       wci_respF_8$ENQ,
       wci_respF_8$FULL_N;

  // ports of submodule wci_respF_9
  reg [33 : 0] wci_respF_9$D_IN;
  wire [33 : 0] wci_respF_9$D_OUT;
  wire wci_respF_9$CLR,
       wci_respF_9$DEQ,
       wci_respF_9$EMPTY_N,
       wci_respF_9$ENQ,
       wci_respF_9$FULL_N;

  // rule scheduling signals
  wire CAN_FIRE_RL_cpDispatch_F_T_F_F,
       CAN_FIRE_RL_cpDispatch_F_T_T_F_F,
       CAN_FIRE_RL_cpDispatch_F_T_T_F_T_F_F,
       CAN_FIRE_RL_cpDispatch_F_T_T_F_T_F_T,
       CAN_FIRE_RL_cpDispatch_F_T_T_F_T_T,
       CAN_FIRE_RL_cpDispatch_F_T_T_T,
       WILL_FIRE_RL_completeWorkerRead,
       WILL_FIRE_RL_completeWorkerWrite,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_T_F,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_T_T,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_F_F_T,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_F_T_F,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_F_T_T,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_T_F,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_T_T,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_F_F_F_T,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_F_F_T,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_F_T_F,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_F_T_T,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_T_F,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_T_T,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_F_F_F_F_T,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_F_F_F_T,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_F_F_T,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_F_T_F,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_F_T_T,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_T_F,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_T_T,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_F_F_F_F_F_F,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_F_F_F_F_F_T,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_F_F_F_F_T,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_F_F_F_T,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_F_F_T,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_F_T_F,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_F_T_T,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_T_F,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_T_T,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_F_F_F_F_F_F,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_F_F_F_F_F_T,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_F_F_F_F_T,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_F_F_F_T,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_F_F_T,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_F_T_F,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_F_T_T,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_T_F,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_T_T,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_F_F_F_F_F_F,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_F_F_F_F_F_T,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_F_F_F_F_T,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_F_F_F_T,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_F_F_T,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_F_T_F,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_F_T_T,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_T_F,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_T_T,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_T_F_F_F_F_F_F,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_T_F_F_F_F_F_T,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_T_F_F_F_F_T,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_T_F_F_F_T,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_T_F_F_T,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_T_F_T_F,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_T_F_T_T,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_T_T_F,
       WILL_FIRE_RL_cpDispatch_F_F_F_F_T_T_T,
       WILL_FIRE_RL_cpDispatch_F_F_F_T,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_F,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_T,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_F,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_F,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_T,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_F,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_F,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_T,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_F,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_F,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_T,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_F,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_T,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_T_F,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_T_T,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_F,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_T,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_F,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_T,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_T_F,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_T_T,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_F_F_F,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_F_F_T,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_F_T_F_F,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_F_T_F_T,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_F_T_T_F,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_T,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_T_F,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_T_T,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_F_F_F,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_F_F_T,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_F_T_F_F,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_F_T_F_T,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_F_T_T_F,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_F_T_T_T,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_T,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_T_F,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_T_T,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_F_F_F,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_F_F_T,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_F_T_F_F,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_F_T_F_T,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_F_T_T_F,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_F_T_T_T,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_T,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_T_F,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_T_T,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_F_F_F,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_F_F_T,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_F_T_F_F,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_F_T_F_T,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_F_T_T_F,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_F_T_T_T,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_T,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_T_F,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_T_T,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_F_F_F,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_F_F_T,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_F_T_F_F,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_F_T_F_T,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_F_T_T_F,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_F_T_T_T,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_T,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_T_F,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_T_T,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_F_F_F_F,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_F_F_F_T,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_F_F_T_F_F,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_F_F_T_F_T,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_F_F_T_T_F,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_F_F_T_T_T,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_F_T,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_T_F,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_T_T,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_F_F_F_F,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_F_F_F_T,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_F_F_T_F_F,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_F_F_T_F_T,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_F_F_T_T_F,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_F_F_T_T_T,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_F_T,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_T_F,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_T_T,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_F_F_F_F,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_F_F_F_T,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_F_F_T_F_F,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_F_F_T_F_T,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_F_F_T_T_F,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_F_F_T_T_T,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_F_T,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_T_F,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_T_T,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_T_F_F_F_F,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_T_F_F_F_T,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_T_F_F_T_F_F,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_T_F_F_T_F_T,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_T_F_F_T_T_F,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_T_F_F_T_T_T,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_T_F_T,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_T_T_F,
       WILL_FIRE_RL_cpDispatch_F_F_T_F_T_T_T,
       WILL_FIRE_RL_cpDispatch_F_F_T_T_F_F_F_F,
       WILL_FIRE_RL_cpDispatch_F_F_T_T_F_F_F_T,
       WILL_FIRE_RL_cpDispatch_F_F_T_T_F_F_T_F_F,
       WILL_FIRE_RL_cpDispatch_F_F_T_T_F_F_T_F_T,
       WILL_FIRE_RL_cpDispatch_F_F_T_T_F_F_T_T_F,
       WILL_FIRE_RL_cpDispatch_F_F_T_T_F_F_T_T_T,
       WILL_FIRE_RL_cpDispatch_F_F_T_T_F_T,
       WILL_FIRE_RL_cpDispatch_F_F_T_T_T_F,
       WILL_FIRE_RL_cpDispatch_F_F_T_T_T_T,
       WILL_FIRE_RL_cpDispatch_F_T_F_T,
       WILL_FIRE_RL_cpDispatch_F_T_T_F_F,
       WILL_FIRE_RL_cpDispatch_F_T_T_F_T_F_F,
       WILL_FIRE_RL_cpDispatch_F_T_T_F_T_F_T,
       WILL_FIRE_RL_cpDispatch_F_T_T_F_T_T,
       WILL_FIRE_RL_cpDispatch_F_T_T_T,
       WILL_FIRE_RL_cpDispatch_T_F_F_F_F_F_F_F_F_F_F,
       WILL_FIRE_RL_cpDispatch_T_F_F_F_F_F_F_F_F_F_T,
       WILL_FIRE_RL_cpDispatch_T_F_F_F_F_F_F_F_F_T,
       WILL_FIRE_RL_cpDispatch_T_F_F_F_F_F_F_F_T,
       WILL_FIRE_RL_cpDispatch_T_F_F_F_F_F_F_T,
       WILL_FIRE_RL_cpDispatch_T_F_F_F_F_F_T,
       WILL_FIRE_RL_cpDispatch_T_F_F_F_F_T_F,
       WILL_FIRE_RL_cpDispatch_T_F_F_F_F_T_T,
       WILL_FIRE_RL_cpDispatch_T_F_F_F_T,
       WILL_FIRE_RL_cpDispatch_T_F_F_T,
       WILL_FIRE_RL_cpDispatch_T_F_T,
       WILL_FIRE_RL_cpDispatch_T_T,
       WILL_FIRE_RL_readAdminResponseCollect,
       WILL_FIRE_RL_reqRcv,
       WILL_FIRE_RL_responseAdminRd,
`ifdef not
       WILL_FIRE_RL_rom_serverAdapter_outData_enqAndDeq,
       WILL_FIRE_RL_rom_serverAdapter_stageReadResponseAlways,
`endif
       WILL_FIRE_RL_wci_reqF_10_both,
       WILL_FIRE_RL_wci_reqF_10_decCtr,
       WILL_FIRE_RL_wci_reqF_10_incCtr,
       WILL_FIRE_RL_wci_reqF_11_both,
       WILL_FIRE_RL_wci_reqF_11_decCtr,
       WILL_FIRE_RL_wci_reqF_11_incCtr,
       WILL_FIRE_RL_wci_reqF_12_both,
       WILL_FIRE_RL_wci_reqF_12_decCtr,
       WILL_FIRE_RL_wci_reqF_12_incCtr,
       WILL_FIRE_RL_wci_reqF_13_both,
       WILL_FIRE_RL_wci_reqF_13_decCtr,
       WILL_FIRE_RL_wci_reqF_13_incCtr,
       WILL_FIRE_RL_wci_reqF_14_both,
       WILL_FIRE_RL_wci_reqF_14_decCtr,
       WILL_FIRE_RL_wci_reqF_14_incCtr,
       WILL_FIRE_RL_wci_reqF_1_both,
       WILL_FIRE_RL_wci_reqF_1_decCtr,
       WILL_FIRE_RL_wci_reqF_1_incCtr,
       WILL_FIRE_RL_wci_reqF_2_both,
       WILL_FIRE_RL_wci_reqF_2_decCtr,
       WILL_FIRE_RL_wci_reqF_2_incCtr,
       WILL_FIRE_RL_wci_reqF_3_both,
       WILL_FIRE_RL_wci_reqF_3_decCtr,
       WILL_FIRE_RL_wci_reqF_3_incCtr,
       WILL_FIRE_RL_wci_reqF_4_both,
       WILL_FIRE_RL_wci_reqF_4_decCtr,
       WILL_FIRE_RL_wci_reqF_4_incCtr,
       WILL_FIRE_RL_wci_reqF_5_both,
       WILL_FIRE_RL_wci_reqF_5_decCtr,
       WILL_FIRE_RL_wci_reqF_5_incCtr,
       WILL_FIRE_RL_wci_reqF_6_both,
       WILL_FIRE_RL_wci_reqF_6_decCtr,
       WILL_FIRE_RL_wci_reqF_6_incCtr,
       WILL_FIRE_RL_wci_reqF_7_both,
       WILL_FIRE_RL_wci_reqF_7_decCtr,
       WILL_FIRE_RL_wci_reqF_7_incCtr,
       WILL_FIRE_RL_wci_reqF_8_both,
       WILL_FIRE_RL_wci_reqF_8_decCtr,
       WILL_FIRE_RL_wci_reqF_8_incCtr,
       WILL_FIRE_RL_wci_reqF_9_both,
       WILL_FIRE_RL_wci_reqF_9_decCtr,
       WILL_FIRE_RL_wci_reqF_9_incCtr,
       WILL_FIRE_RL_wci_reqF_both,
       WILL_FIRE_RL_wci_reqF_decCtr,
       WILL_FIRE_RL_wci_reqF_incCtr,
       WILL_FIRE_RL_wci_wrkBusy,
       WILL_FIRE_RL_wci_wrkBusy_1,
       WILL_FIRE_RL_wci_wrkBusy_10,
       WILL_FIRE_RL_wci_wrkBusy_11,
       WILL_FIRE_RL_wci_wrkBusy_12,
       WILL_FIRE_RL_wci_wrkBusy_13,
       WILL_FIRE_RL_wci_wrkBusy_14,
       WILL_FIRE_RL_wci_wrkBusy_2,
       WILL_FIRE_RL_wci_wrkBusy_3,
       WILL_FIRE_RL_wci_wrkBusy_4,
       WILL_FIRE_RL_wci_wrkBusy_5,
       WILL_FIRE_RL_wci_wrkBusy_6,
       WILL_FIRE_RL_wci_wrkBusy_7,
       WILL_FIRE_RL_wci_wrkBusy_8,
       WILL_FIRE_RL_wci_wrkBusy_9;

  // inputs to muxes for submodule ports
  reg [71 : 0] MUX_wci_reqF_10_q_0$write_1__VAL_1,
	       MUX_wci_reqF_11_q_0$write_1__VAL_1,
	       MUX_wci_reqF_12_q_0$write_1__VAL_1,
	       MUX_wci_reqF_13_q_0$write_1__VAL_1,
	       MUX_wci_reqF_14_q_0$write_1__VAL_1,
	       MUX_wci_reqF_1_q_0$write_1__VAL_2,
	       MUX_wci_reqF_2_q_0$write_1__VAL_2,
	       MUX_wci_reqF_3_q_0$write_1__VAL_2,
	       MUX_wci_reqF_4_q_0$write_1__VAL_2,
	       MUX_wci_reqF_5_q_0$write_1__VAL_2,
	       MUX_wci_reqF_6_q_0$write_1__VAL_2,
	       MUX_wci_reqF_7_q_0$write_1__VAL_2,
	       MUX_wci_reqF_8_q_0$write_1__VAL_2,
	       MUX_wci_reqF_9_q_0$write_1__VAL_2,
	       MUX_wci_reqF_q_0$write_1__VAL_2;
  reg [2 : 0] MUX_wci_reqERR$write_1__VAL_1,
	      MUX_wci_reqERR_1$write_1__VAL_1,
	      MUX_wci_reqERR_10$write_1__VAL_1,
	      MUX_wci_reqERR_11$write_1__VAL_1,
	      MUX_wci_reqERR_12$write_1__VAL_1,
	      MUX_wci_reqERR_13$write_1__VAL_1,
	      MUX_wci_reqERR_14$write_1__VAL_1,
	      MUX_wci_reqERR_2$write_1__VAL_1,
	      MUX_wci_reqERR_3$write_1__VAL_1,
	      MUX_wci_reqERR_4$write_1__VAL_1,
	      MUX_wci_reqERR_5$write_1__VAL_1,
	      MUX_wci_reqERR_6$write_1__VAL_1,
	      MUX_wci_reqERR_7$write_1__VAL_1,
	      MUX_wci_reqERR_8$write_1__VAL_1,
	      MUX_wci_reqERR_9$write_1__VAL_1,
	      MUX_wci_reqFAIL$write_1__VAL_1,
	      MUX_wci_reqFAIL_1$write_1__VAL_1,
	      MUX_wci_reqFAIL_10$write_1__VAL_1,
	      MUX_wci_reqFAIL_11$write_1__VAL_1,
	      MUX_wci_reqFAIL_12$write_1__VAL_1,
	      MUX_wci_reqFAIL_13$write_1__VAL_1,
	      MUX_wci_reqFAIL_14$write_1__VAL_1,
	      MUX_wci_reqFAIL_2$write_1__VAL_1,
	      MUX_wci_reqFAIL_3$write_1__VAL_1,
	      MUX_wci_reqFAIL_4$write_1__VAL_1,
	      MUX_wci_reqFAIL_5$write_1__VAL_1,
	      MUX_wci_reqFAIL_6$write_1__VAL_1,
	      MUX_wci_reqFAIL_7$write_1__VAL_1,
	      MUX_wci_reqFAIL_8$write_1__VAL_1,
	      MUX_wci_reqFAIL_9$write_1__VAL_1,
	      MUX_wci_reqTO$write_1__VAL_1,
	      MUX_wci_reqTO_1$write_1__VAL_1,
	      MUX_wci_reqTO_10$write_1__VAL_1,
	      MUX_wci_reqTO_11$write_1__VAL_1,
	      MUX_wci_reqTO_12$write_1__VAL_1,
	      MUX_wci_reqTO_13$write_1__VAL_1,
	      MUX_wci_reqTO_14$write_1__VAL_1,
	      MUX_wci_reqTO_2$write_1__VAL_1,
	      MUX_wci_reqTO_3$write_1__VAL_1,
	      MUX_wci_reqTO_4$write_1__VAL_1,
	      MUX_wci_reqTO_5$write_1__VAL_1,
	      MUX_wci_reqTO_6$write_1__VAL_1,
	      MUX_wci_reqTO_7$write_1__VAL_1,
	      MUX_wci_reqTO_8$write_1__VAL_1,
	      MUX_wci_reqTO_9$write_1__VAL_1;
  wire [71 : 0] MUX_wci_reqF_10_q_0$write_1__VAL_2,
		MUX_wci_reqF_10_x_wire$wset_1__VAL_1,
		MUX_wci_reqF_10_x_wire$wset_1__VAL_2,
		MUX_wci_reqF_10_x_wire$wset_1__VAL_3,
		MUX_wci_reqF_11_q_0$write_1__VAL_2,
		MUX_wci_reqF_11_x_wire$wset_1__VAL_1,
		MUX_wci_reqF_11_x_wire$wset_1__VAL_2,
		MUX_wci_reqF_12_q_0$write_1__VAL_2,
		MUX_wci_reqF_12_x_wire$wset_1__VAL_1,
		MUX_wci_reqF_12_x_wire$wset_1__VAL_2,
		MUX_wci_reqF_13_q_0$write_1__VAL_2,
		MUX_wci_reqF_13_x_wire$wset_1__VAL_1,
		MUX_wci_reqF_13_x_wire$wset_1__VAL_2,
		MUX_wci_reqF_14_q_0$write_1__VAL_2,
		MUX_wci_reqF_14_x_wire$wset_1__VAL_1,
		MUX_wci_reqF_14_x_wire$wset_1__VAL_2,
		MUX_wci_reqF_1_q_0$write_1__VAL_1,
		MUX_wci_reqF_1_x_wire$wset_1__VAL_1,
		MUX_wci_reqF_1_x_wire$wset_1__VAL_2,
		MUX_wci_reqF_2_q_0$write_1__VAL_1,
		MUX_wci_reqF_2_x_wire$wset_1__VAL_1,
		MUX_wci_reqF_2_x_wire$wset_1__VAL_2,
		MUX_wci_reqF_3_q_0$write_1__VAL_1,
		MUX_wci_reqF_3_x_wire$wset_1__VAL_1,
		MUX_wci_reqF_3_x_wire$wset_1__VAL_2,
		MUX_wci_reqF_4_q_0$write_1__VAL_1,
		MUX_wci_reqF_4_x_wire$wset_1__VAL_1,
		MUX_wci_reqF_4_x_wire$wset_1__VAL_2,
		MUX_wci_reqF_5_q_0$write_1__VAL_1,
		MUX_wci_reqF_5_x_wire$wset_1__VAL_1,
		MUX_wci_reqF_5_x_wire$wset_1__VAL_2,
		MUX_wci_reqF_6_q_0$write_1__VAL_1,
		MUX_wci_reqF_6_x_wire$wset_1__VAL_1,
		MUX_wci_reqF_6_x_wire$wset_1__VAL_2,
		MUX_wci_reqF_7_q_0$write_1__VAL_1,
		MUX_wci_reqF_7_x_wire$wset_1__VAL_1,
		MUX_wci_reqF_7_x_wire$wset_1__VAL_2,
		MUX_wci_reqF_8_q_0$write_1__VAL_1,
		MUX_wci_reqF_8_x_wire$wset_1__VAL_1,
		MUX_wci_reqF_8_x_wire$wset_1__VAL_2,
		MUX_wci_reqF_9_q_0$write_1__VAL_1,
		MUX_wci_reqF_9_x_wire$wset_1__VAL_1,
		MUX_wci_reqF_9_x_wire$wset_1__VAL_2,
		MUX_wci_reqF_q_0$write_1__VAL_1,
		MUX_wci_reqF_x_wire$wset_1__VAL_1,
		MUX_wci_reqF_x_wire$wset_1__VAL_2;
  wire [64 : 0] MUX_cpReq$write_1__VAL_4;
  wire [39 : 0] MUX_cpRespF$enq_1__VAL_1, MUX_cpRespF$enq_1__VAL_2;
  wire [33 : 0] MUX_wci_respF$enq_1__VAL_1,
		MUX_wci_respF$enq_1__VAL_2,
		MUX_wci_respF$enq_1__VAL_3,
		MUX_wci_respF$enq_1__VAL_4,
		MUX_wci_respF$enq_1__VAL_5,
		MUX_wci_respF_1$enq_1__VAL_1,
		MUX_wci_respF_1$enq_1__VAL_2,
		MUX_wci_respF_1$enq_1__VAL_3,
		MUX_wci_respF_1$enq_1__VAL_4,
		MUX_wci_respF_1$enq_1__VAL_5,
		MUX_wci_respF_10$enq_1__VAL_1,
		MUX_wci_respF_10$enq_1__VAL_2,
		MUX_wci_respF_10$enq_1__VAL_3,
		MUX_wci_respF_10$enq_1__VAL_4,
		MUX_wci_respF_10$enq_1__VAL_5,
		MUX_wci_respF_11$enq_1__VAL_1,
		MUX_wci_respF_11$enq_1__VAL_2,
		MUX_wci_respF_11$enq_1__VAL_3,
		MUX_wci_respF_11$enq_1__VAL_4,
		MUX_wci_respF_11$enq_1__VAL_5,
		MUX_wci_respF_12$enq_1__VAL_1,
		MUX_wci_respF_12$enq_1__VAL_2,
		MUX_wci_respF_12$enq_1__VAL_3,
		MUX_wci_respF_12$enq_1__VAL_4,
		MUX_wci_respF_12$enq_1__VAL_5,
		MUX_wci_respF_13$enq_1__VAL_1,
		MUX_wci_respF_13$enq_1__VAL_2,
		MUX_wci_respF_13$enq_1__VAL_3,
		MUX_wci_respF_13$enq_1__VAL_4,
		MUX_wci_respF_13$enq_1__VAL_5,
		MUX_wci_respF_14$enq_1__VAL_1,
		MUX_wci_respF_14$enq_1__VAL_2,
		MUX_wci_respF_14$enq_1__VAL_3,
		MUX_wci_respF_14$enq_1__VAL_4,
		MUX_wci_respF_14$enq_1__VAL_5,
		MUX_wci_respF_2$enq_1__VAL_1,
		MUX_wci_respF_2$enq_1__VAL_2,
		MUX_wci_respF_2$enq_1__VAL_3,
		MUX_wci_respF_2$enq_1__VAL_4,
		MUX_wci_respF_2$enq_1__VAL_5,
		MUX_wci_respF_3$enq_1__VAL_1,
		MUX_wci_respF_3$enq_1__VAL_2,
		MUX_wci_respF_3$enq_1__VAL_3,
		MUX_wci_respF_3$enq_1__VAL_4,
		MUX_wci_respF_3$enq_1__VAL_5,
		MUX_wci_respF_4$enq_1__VAL_1,
		MUX_wci_respF_4$enq_1__VAL_2,
		MUX_wci_respF_4$enq_1__VAL_3,
		MUX_wci_respF_4$enq_1__VAL_4,
		MUX_wci_respF_4$enq_1__VAL_5,
		MUX_wci_respF_5$enq_1__VAL_1,
		MUX_wci_respF_5$enq_1__VAL_2,
		MUX_wci_respF_5$enq_1__VAL_3,
		MUX_wci_respF_5$enq_1__VAL_4,
		MUX_wci_respF_5$enq_1__VAL_5,
		MUX_wci_respF_6$enq_1__VAL_1,
		MUX_wci_respF_6$enq_1__VAL_2,
		MUX_wci_respF_6$enq_1__VAL_3,
		MUX_wci_respF_6$enq_1__VAL_4,
		MUX_wci_respF_6$enq_1__VAL_5,
		MUX_wci_respF_7$enq_1__VAL_1,
		MUX_wci_respF_7$enq_1__VAL_2,
		MUX_wci_respF_7$enq_1__VAL_3,
		MUX_wci_respF_7$enq_1__VAL_4,
		MUX_wci_respF_7$enq_1__VAL_5,
		MUX_wci_respF_8$enq_1__VAL_1,
		MUX_wci_respF_8$enq_1__VAL_2,
		MUX_wci_respF_8$enq_1__VAL_3,
		MUX_wci_respF_8$enq_1__VAL_4,
		MUX_wci_respF_8$enq_1__VAL_5,
		MUX_wci_respF_9$enq_1__VAL_1,
		MUX_wci_respF_9$enq_1__VAL_2,
		MUX_wci_respF_9$enq_1__VAL_3,
		MUX_wci_respF_9$enq_1__VAL_4,
		MUX_wci_respF_9$enq_1__VAL_5;
  wire [32 : 0] MUX_adminResp2F$enq_1__VAL_1,
		MUX_adminResp2F$enq_1__VAL_2,
		MUX_adminResp2F$enq_1__VAL_3;
  wire [31 : 0] MUX_readCntReg$write_1__VAL_2,
		MUX_wci_respTimr$write_1__VAL_2,
		MUX_wci_respTimr_1$write_1__VAL_2,
		MUX_wci_respTimr_10$write_1__VAL_2,
		MUX_wci_respTimr_11$write_1__VAL_2,
		MUX_wci_respTimr_12$write_1__VAL_2,
		MUX_wci_respTimr_13$write_1__VAL_2,
		MUX_wci_respTimr_14$write_1__VAL_2,
		MUX_wci_respTimr_2$write_1__VAL_2,
		MUX_wci_respTimr_3$write_1__VAL_2,
		MUX_wci_respTimr_4$write_1__VAL_2,
		MUX_wci_respTimr_5$write_1__VAL_2,
		MUX_wci_respTimr_6$write_1__VAL_2,
		MUX_wci_respTimr_7$write_1__VAL_2,
		MUX_wci_respTimr_8$write_1__VAL_2,
		MUX_wci_respTimr_9$write_1__VAL_2;
  wire MUX_wci_busy$write_1__SEL_1,
       MUX_wci_busy$write_1__SEL_2,
       MUX_wci_busy_1$write_1__SEL_1,
       MUX_wci_busy_1$write_1__SEL_2,
       MUX_wci_busy_10$write_1__SEL_1,
       MUX_wci_busy_10$write_1__SEL_2,
       MUX_wci_busy_11$write_1__SEL_1,
       MUX_wci_busy_11$write_1__SEL_2,
       MUX_wci_busy_12$write_1__SEL_1,
       MUX_wci_busy_12$write_1__SEL_2,
       MUX_wci_busy_13$write_1__SEL_1,
       MUX_wci_busy_13$write_1__SEL_2,
       MUX_wci_busy_14$write_1__SEL_1,
       MUX_wci_busy_14$write_1__SEL_2,
       MUX_wci_busy_2$write_1__SEL_1,
       MUX_wci_busy_2$write_1__SEL_2,
       MUX_wci_busy_3$write_1__SEL_1,
       MUX_wci_busy_3$write_1__SEL_2,
       MUX_wci_busy_4$write_1__SEL_1,
       MUX_wci_busy_4$write_1__SEL_2,
       MUX_wci_busy_5$write_1__SEL_1,
       MUX_wci_busy_5$write_1__SEL_2,
       MUX_wci_busy_6$write_1__SEL_1,
       MUX_wci_busy_6$write_1__SEL_2,
       MUX_wci_busy_7$write_1__SEL_1,
       MUX_wci_busy_7$write_1__SEL_2,
       MUX_wci_busy_8$write_1__SEL_1,
       MUX_wci_busy_8$write_1__SEL_2,
       MUX_wci_busy_9$write_1__SEL_1,
       MUX_wci_busy_9$write_1__SEL_2,
       MUX_wci_reqERR$write_1__SEL_1,
       MUX_wci_reqERR_1$write_1__SEL_1,
       MUX_wci_reqERR_10$write_1__SEL_1,
       MUX_wci_reqERR_11$write_1__SEL_1,
       MUX_wci_reqERR_12$write_1__SEL_1,
       MUX_wci_reqERR_13$write_1__SEL_1,
       MUX_wci_reqERR_14$write_1__SEL_1,
       MUX_wci_reqERR_2$write_1__SEL_1,
       MUX_wci_reqERR_3$write_1__SEL_1,
       MUX_wci_reqERR_4$write_1__SEL_1,
       MUX_wci_reqERR_5$write_1__SEL_1,
       MUX_wci_reqERR_6$write_1__SEL_1,
       MUX_wci_reqERR_7$write_1__SEL_1,
       MUX_wci_reqERR_8$write_1__SEL_1,
       MUX_wci_reqERR_9$write_1__SEL_1,
       MUX_wci_reqFAIL$write_1__SEL_1,
       MUX_wci_reqFAIL_1$write_1__SEL_1,
       MUX_wci_reqFAIL_10$write_1__SEL_1,
       MUX_wci_reqFAIL_11$write_1__SEL_1,
       MUX_wci_reqFAIL_12$write_1__SEL_1,
       MUX_wci_reqFAIL_13$write_1__SEL_1,
       MUX_wci_reqFAIL_14$write_1__SEL_1,
       MUX_wci_reqFAIL_2$write_1__SEL_1,
       MUX_wci_reqFAIL_3$write_1__SEL_1,
       MUX_wci_reqFAIL_4$write_1__SEL_1,
       MUX_wci_reqFAIL_5$write_1__SEL_1,
       MUX_wci_reqFAIL_6$write_1__SEL_1,
       MUX_wci_reqFAIL_7$write_1__SEL_1,
       MUX_wci_reqFAIL_8$write_1__SEL_1,
       MUX_wci_reqFAIL_9$write_1__SEL_1,
       MUX_wci_reqF_10_c_r$write_1__VAL_1,
       MUX_wci_reqF_10_c_r$write_1__VAL_2,
       MUX_wci_reqF_10_q_0$write_1__SEL_1,
       MUX_wci_reqF_11_c_r$write_1__VAL_1,
       MUX_wci_reqF_11_c_r$write_1__VAL_2,
       MUX_wci_reqF_11_q_0$write_1__SEL_1,
       MUX_wci_reqF_12_c_r$write_1__VAL_1,
       MUX_wci_reqF_12_c_r$write_1__VAL_2,
       MUX_wci_reqF_12_q_0$write_1__SEL_1,
       MUX_wci_reqF_13_c_r$write_1__VAL_1,
       MUX_wci_reqF_13_c_r$write_1__VAL_2,
       MUX_wci_reqF_13_q_0$write_1__SEL_1,
       MUX_wci_reqF_14_c_r$write_1__VAL_1,
       MUX_wci_reqF_14_c_r$write_1__VAL_2,
       MUX_wci_reqF_14_q_0$write_1__SEL_1,
       MUX_wci_reqF_1_c_r$write_1__VAL_1,
       MUX_wci_reqF_1_c_r$write_1__VAL_2,
       MUX_wci_reqF_1_q_0$write_1__SEL_2,
       MUX_wci_reqF_2_c_r$write_1__VAL_1,
       MUX_wci_reqF_2_c_r$write_1__VAL_2,
       MUX_wci_reqF_2_q_0$write_1__SEL_2,
       MUX_wci_reqF_3_c_r$write_1__VAL_1,
       MUX_wci_reqF_3_c_r$write_1__VAL_2,
       MUX_wci_reqF_3_q_0$write_1__SEL_2,
       MUX_wci_reqF_4_c_r$write_1__VAL_1,
       MUX_wci_reqF_4_c_r$write_1__VAL_2,
       MUX_wci_reqF_4_q_0$write_1__SEL_2,
       MUX_wci_reqF_5_c_r$write_1__VAL_1,
       MUX_wci_reqF_5_c_r$write_1__VAL_2,
       MUX_wci_reqF_5_q_0$write_1__SEL_2,
       MUX_wci_reqF_6_c_r$write_1__VAL_1,
       MUX_wci_reqF_6_c_r$write_1__VAL_2,
       MUX_wci_reqF_6_q_0$write_1__SEL_2,
       MUX_wci_reqF_7_c_r$write_1__VAL_1,
       MUX_wci_reqF_7_c_r$write_1__VAL_2,
       MUX_wci_reqF_7_q_0$write_1__SEL_2,
       MUX_wci_reqF_8_c_r$write_1__VAL_1,
       MUX_wci_reqF_8_c_r$write_1__VAL_2,
       MUX_wci_reqF_8_q_0$write_1__SEL_2,
       MUX_wci_reqF_9_c_r$write_1__VAL_1,
       MUX_wci_reqF_9_c_r$write_1__VAL_2,
       MUX_wci_reqF_9_q_0$write_1__SEL_2,
       MUX_wci_reqF_c_r$write_1__VAL_1,
       MUX_wci_reqF_c_r$write_1__VAL_2,
       MUX_wci_reqF_q_0$write_1__SEL_2,
       MUX_wci_reqPend$write_1__SEL_1,
       MUX_wci_reqPend_1$write_1__SEL_1,
       MUX_wci_reqPend_10$write_1__SEL_1,
       MUX_wci_reqPend_11$write_1__SEL_1,
       MUX_wci_reqPend_12$write_1__SEL_1,
       MUX_wci_reqPend_13$write_1__SEL_1,
       MUX_wci_reqPend_14$write_1__SEL_1,
       MUX_wci_reqPend_2$write_1__SEL_1,
       MUX_wci_reqPend_3$write_1__SEL_1,
       MUX_wci_reqPend_4$write_1__SEL_1,
       MUX_wci_reqPend_5$write_1__SEL_1,
       MUX_wci_reqPend_6$write_1__SEL_1,
       MUX_wci_reqPend_7$write_1__SEL_1,
       MUX_wci_reqPend_8$write_1__SEL_1,
       MUX_wci_reqPend_9$write_1__SEL_1,
       MUX_wci_reqTO$write_1__SEL_1,
       MUX_wci_reqTO_1$write_1__SEL_1,
       MUX_wci_reqTO_10$write_1__SEL_1,
       MUX_wci_reqTO_11$write_1__SEL_1,
       MUX_wci_reqTO_12$write_1__SEL_1,
       MUX_wci_reqTO_13$write_1__SEL_1,
       MUX_wci_reqTO_14$write_1__SEL_1,
       MUX_wci_reqTO_2$write_1__SEL_1,
       MUX_wci_reqTO_3$write_1__SEL_1,
       MUX_wci_reqTO_4$write_1__SEL_1,
       MUX_wci_reqTO_5$write_1__SEL_1,
       MUX_wci_reqTO_6$write_1__SEL_1,
       MUX_wci_reqTO_7$write_1__SEL_1,
       MUX_wci_reqTO_8$write_1__SEL_1,
       MUX_wci_reqTO_9$write_1__SEL_1,
       MUX_wci_respF$enq_1__SEL_6,
       MUX_wci_respF$enq_1__SEL_7,
       MUX_wci_respF_1$enq_1__SEL_6,
       MUX_wci_respF_1$enq_1__SEL_7,
       MUX_wci_respF_10$enq_1__SEL_6,
       MUX_wci_respF_10$enq_1__SEL_7,
       MUX_wci_respF_11$enq_1__SEL_6,
       MUX_wci_respF_11$enq_1__SEL_7,
       MUX_wci_respF_12$enq_1__SEL_6,
       MUX_wci_respF_12$enq_1__SEL_7,
       MUX_wci_respF_13$enq_1__SEL_6,
       MUX_wci_respF_13$enq_1__SEL_7,
       MUX_wci_respF_14$enq_1__SEL_6,
       MUX_wci_respF_14$enq_1__SEL_7,
       MUX_wci_respF_2$enq_1__SEL_6,
       MUX_wci_respF_2$enq_1__SEL_7,
       MUX_wci_respF_3$enq_1__SEL_6,
       MUX_wci_respF_3$enq_1__SEL_7,
       MUX_wci_respF_4$enq_1__SEL_6,
       MUX_wci_respF_4$enq_1__SEL_7,
       MUX_wci_respF_5$enq_1__SEL_6,
       MUX_wci_respF_5$enq_1__SEL_7,
       MUX_wci_respF_6$enq_1__SEL_6,
       MUX_wci_respF_6$enq_1__SEL_7,
       MUX_wci_respF_7$enq_1__SEL_6,
       MUX_wci_respF_7$enq_1__SEL_7,
       MUX_wci_respF_8$enq_1__SEL_6,
       MUX_wci_respF_8$enq_1__SEL_7,
       MUX_wci_respF_9$enq_1__SEL_6,
       MUX_wci_respF_9$enq_1__SEL_7,
       MUX_wrkAct$write_1__SEL_1,
       MUX_wrkAct$write_1__SEL_2,
       MUX_wrkAct$write_1__SEL_3;

  // remaining internal signals
  reg [63 : 0] v__h106118,
	       v__h106171,
	       v__h12057,
	       v__h12147,
	       v__h12236,
	       v__h12460,
	       v__h12550,
	       v__h12639,
	       v__h12868,
	       v__h12958,
	       v__h13047,
	       v__h16497,
	       v__h16587,
	       v__h16676,
	       v__h16900,
	       v__h16990,
	       v__h17079,
	       v__h17308,
	       v__h17398,
	       v__h17487,
	       v__h20937,
	       v__h21027,
	       v__h21116,
	       v__h21340,
	       v__h21430,
	       v__h21519,
	       v__h21748,
	       v__h21838,
	       v__h21927,
	       v__h25377,
	       v__h25467,
	       v__h25556,
	       v__h25780,
	       v__h25870,
	       v__h25959,
	       v__h26188,
	       v__h26278,
	       v__h26367,
	       v__h29817,
	       v__h29907,
	       v__h29996,
	       v__h30220,
	       v__h30310,
	       v__h30399,
	       v__h30628,
	       v__h30718,
	       v__h30807,
	       v__h34257,
	       v__h34347,
	       v__h34436,
	       v__h34660,
	       v__h34750,
	       v__h34839,
	       v__h35068,
	       v__h35158,
	       v__h35247,
	       v__h38697,
	       v__h38787,
	       v__h38876,
	       v__h39100,
	       v__h39190,
	       v__h39279,
	       v__h39508,
	       v__h39598,
	       v__h39687,
	       v__h43137,
	       v__h43227,
	       v__h43316,
	       v__h43540,
	       v__h43630,
	       v__h43719,
	       v__h43948,
	       v__h44038,
	       v__h44127,
	       v__h47577,
	       v__h47667,
	       v__h47756,
	       v__h47980,
	       v__h48070,
	       v__h48159,
	       v__h48388,
	       v__h48478,
	       v__h48567,
	       v__h52017,
	       v__h52107,
	       v__h52196,
	       v__h52420,
	       v__h52510,
	       v__h52599,
	       v__h52828,
	       v__h52918,
	       v__h53007,
	       v__h56457,
	       v__h56547,
	       v__h56636,
	       v__h56860,
	       v__h56950,
	       v__h57039,
	       v__h57268,
	       v__h57358,
	       v__h57447,
	       v__h60897,
	       v__h60987,
	       v__h61076,
	       v__h61300,
	       v__h61390,
	       v__h61479,
	       v__h61708,
	       v__h61798,
	       v__h61887,
	       v__h65337,
	       v__h65427,
	       v__h65516,
	       v__h65740,
	       v__h65830,
	       v__h65919,
	       v__h66148,
	       v__h66238,
	       v__h66327,
	       v__h69777,
	       v__h69867,
	       v__h69956,
	       v__h70180,
	       v__h70270,
	       v__h70359,
	       v__h70588,
	       v__h70678,
	       v__h70767,
	       v__h74217,
	       v__h74307,
	       v__h74396,
	       v__h74620,
	       v__h74710,
	       v__h74799,
	       v__h75028,
	       v__h75118,
	       v__h75207,
	       v__h79502,
	       v__h80094,
	       v__h80203,
	       v__h80782,
	       v__h80891,
	       v__h81470,
	       v__h81579,
	       v__h82158,
	       v__h82267,
	       v__h82846,
	       v__h82955,
	       v__h83534,
	       v__h83643,
	       v__h84222,
	       v__h84331,
	       v__h84910,
	       v__h85019,
	       v__h85598,
	       v__h85707,
	       v__h86286,
	       v__h86395,
	       v__h86974,
	       v__h87083,
	       v__h87662,
	       v__h87771,
	       v__h88350,
	       v__h88459,
	       v__h89038,
	       v__h89147,
	       v__h89726,
	       v__h97130,
	       v__h97202,
	       v__h97274,
	       v__h97346,
	       v__h97418,
	       v__h97490,
	       v__h97562,
	       v__h97634,
	       v__h97706,
	       v__h97778,
	       v__h97850,
	       v__h97922,
	       v__h97994,
	       v__h98066,
	       v__h98138;
  reg [31 : 0] CASE_cpReq_BITS_9_TO_6_uuid_arg_BITS_31_TO_0_0_ETC__q3,
	       IF_cpReq_363_BITS_11_TO_4_366_EQ_0x0_445_THEN__ETC___d6178,
	       IF_cpReq_363_BITS_11_TO_4_366_EQ_0x30_595_THEN_ETC___d6177,
	       rtnData__h113334;
  reg IF_wrkAct_077_EQ_0_078_THEN_wci_respF_i_notEmp_ETC___d6132;
`ifdef not
  wire [49 : 0] _281474976710656_MINUS_timeServ_delSecond__q1,
		x__h3700,
		x__h4421,
		x__h4649;
`endif
  wire [47 : 0] x_f__h4848;
  wire [32 : 0] IF_adminResp2F_notEmpty__304_THEN_adminResp2F__ETC___d2342;
  wire [31 : 0] cpStatus__h75932,
		crr_data__h76602,
		toCount__h11764,
		toCount__h16210,
		toCount__h20650,
		toCount__h25090,
		toCount__h29530,
		toCount__h33970,
		toCount__h38410,
		toCount__h42850,
		toCount__h47290,
		toCount__h51730,
		toCount__h56170,
		toCount__h60610,
		toCount__h65050,
		toCount__h69490,
		toCount__h73930,
		wciAddr__h78327,
		wciAddr__h78395,
		wciAddr__h78461,
		wciAddr__h78527,
		wciAddr__h78593,
		wciAddr__h78659,
		wciAddr__h78725,
		wciAddr__h78791,
		wciAddr__h78857,
		wciAddr__h78923,
		wciAddr__h78989,
		wciAddr__h79055,
		wciAddr__h79121,
		wciAddr__h79187,
		wciAddr__h79253,
		x__h11924,
		x__h16367,
		x__h20807,
		x__h25247,
		x__h29687,
		x__h34127,
		x__h38567,
		x__h43007,
`ifdef not
		x__h4715,
`endif
		x__h47447,
		x__h51887,
		x__h56327,
		x__h60767,
		x__h65207,
		x__h69647,
		x__h74087,
		x_addr__h98551,
		x_data__h104757,
		x_data__h104763,
		x_data__h104810,
		x_data__h104816,
		x_data__h104863,
		x_data__h104869,
		x_data__h104916,
		x_data__h104922,
		x_data__h104969,
		x_data__h104975,
		x_data__h105022,
		x_data__h105028,
		x_data__h105075,
		x_data__h105081,
		x_data__h105128,
		x_data__h105134,
		x_data__h105181,
		x_data__h105187,
		x_data__h105234,
		x_data__h105240,
		x_data__h105287,
		x_data__h105293,
		x_data__h105340,
		x_data__h105346,
		x_data__h105393,
		x_data__h105399,
		x_data__h105446,
		x_data__h105452,
		x_data__h105499,
		x_data__h105505;
  wire [26 : 0] IF_wci_lastControlOp_10_713_BIT_3_714_THEN_wci_ETC___d1728,
		IF_wci_lastControlOp_11_853_BIT_3_854_THEN_wci_ETC___d1868,
		IF_wci_lastControlOp_12_993_BIT_3_994_THEN_wci_ETC___d2008,
		IF_wci_lastControlOp_13_133_BIT_3_134_THEN_wci_ETC___d2148,
		IF_wci_lastControlOp_13_BIT_3_14_THEN_wci_last_ETC___d328,
		IF_wci_lastControlOp_14_273_BIT_3_274_THEN_wci_ETC___d2288,
		IF_wci_lastControlOp_1_53_BIT_3_54_THEN_wci_la_ETC___d468,
		IF_wci_lastControlOp_2_93_BIT_3_94_THEN_wci_la_ETC___d608,
		IF_wci_lastControlOp_3_33_BIT_3_34_THEN_wci_la_ETC___d748,
		IF_wci_lastControlOp_4_73_BIT_3_74_THEN_wci_la_ETC___d888,
		IF_wci_lastControlOp_5_013_BIT_3_014_THEN_wci__ETC___d1028,
		IF_wci_lastControlOp_6_153_BIT_3_154_THEN_wci__ETC___d1168,
		IF_wci_lastControlOp_7_293_BIT_3_294_THEN_wci__ETC___d1308,
		IF_wci_lastControlOp_8_433_BIT_3_434_THEN_wci__ETC___d1448,
		IF_wci_lastControlOp_9_573_BIT_3_574_THEN_wci__ETC___d1588;
  wire [23 : 0] bAddr__h113843, bAddr__h114303;
`ifdef not
  wire [21 : 0] _281474976710656_MINUS_timeServ_delSecond_BITS__ETC__q2;
`endif
  wire [14 : 0] x__h106341, x__h106890;
  wire [4 : 0] x__h98553;
  wire [3 : 0] _theResult_____1__h76796,
	       _theResult_____1__h76814,
	       wn___1__h77585,
	       wn__h76795;
`ifdef not
  wire [2 : 0] rom_serverAdapter_cnt_29_PLUS_IF_rom_serverAda_ETC___d135;
`endif
  wire IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d3932,
       IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d3941,
       IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d3951,
       IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4010,
       IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4019,
       IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4029,
       IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4086,
       IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4095,
       IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4105,
       IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4162,
       IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4171,
       IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4181,
       IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4238,
       IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4247,
       IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4257,
       IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4314,
       IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4323,
       IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4333,
       IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4390,
       IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4399,
       IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4409,
       IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4466,
       IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4475,
       IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4485,
       IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4542,
       IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4551,
       IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4561,
       IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4618,
       IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4627,
       IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4637,
       IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4694,
       IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4703,
       IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4713,
       IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4770,
       IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4779,
       IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4789,
       IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4846,
       IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4855,
       IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4865,
       IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4922,
       IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4931,
       IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4941,
       IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4998,
       IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d5007,
       IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d5017,
`ifdef not
       IF_timeServ_ppsOK_7_THEN_timeServ_ppsExtSync_d_ETC___d5465,
`endif
       NOT_cpReq_363_BITS_11_TO_4_366_EQ_0x30_595_649_ETC___d2712,
       NOT_cpReq_363_BITS_64_TO_62_364_EQ_0_881_886_A_ETC___d5073,
       NOT_cpReq_363_BITS_64_TO_62_364_EQ_3_877_885_A_ETC___d3976,
       NOT_cpReq_363_BITS_64_TO_62_364_EQ_3_877_885_A_ETC___d4052,
       NOT_cpReq_363_BITS_64_TO_62_364_EQ_3_877_885_A_ETC___d4128,
       NOT_cpReq_363_BITS_64_TO_62_364_EQ_3_877_885_A_ETC___d4204,
       NOT_cpReq_363_BITS_64_TO_62_364_EQ_3_877_885_A_ETC___d4280,
       NOT_cpReq_363_BITS_64_TO_62_364_EQ_3_877_885_A_ETC___d4356,
       NOT_cpReq_363_BITS_64_TO_62_364_EQ_3_877_885_A_ETC___d4432,
       NOT_cpReq_363_BITS_64_TO_62_364_EQ_3_877_885_A_ETC___d4508,
       NOT_cpReq_363_BITS_64_TO_62_364_EQ_3_877_885_A_ETC___d4584,
       NOT_cpReq_363_BITS_64_TO_62_364_EQ_3_877_885_A_ETC___d4660,
       NOT_cpReq_363_BITS_64_TO_62_364_EQ_3_877_885_A_ETC___d4736,
       NOT_cpReq_363_BITS_64_TO_62_364_EQ_3_877_885_A_ETC___d4812,
       NOT_cpReq_363_BITS_64_TO_62_364_EQ_3_877_885_A_ETC___d4888,
       NOT_cpReq_363_BITS_64_TO_62_364_EQ_3_877_885_A_ETC___d4964,
       NOT_cpReq_363_BITS_64_TO_62_364_EQ_3_877_885_A_ETC___d5040,
       NOT_cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_961_A_ETC___d2962,
       NOT_cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_961_A_ETC___d3025,
       NOT_cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_961_A_ETC___d3088,
       NOT_cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_961_A_ETC___d3151,
       NOT_cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_961_A_ETC___d3214,
       NOT_cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_961_A_ETC___d3277,
       NOT_cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_961_A_ETC___d3340,
       NOT_cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_961_A_ETC___d3403,
       NOT_cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_961_A_ETC___d3466,
       NOT_cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_961_A_ETC___d3529,
       NOT_cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_961_A_ETC___d3592,
       NOT_cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_961_A_ETC___d3655,
       NOT_cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_961_A_ETC___d3718,
       NOT_cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_961_A_ETC___d3781,
       NOT_cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_961_A_ETC___d3844,
       NOT_cpReq_363_BIT_36_924_932_AND_NOT_wci_busy__ETC___d2933,
       NOT_cpReq_363_BIT_36_924_932_AND_NOT_wci_busy__ETC___d3000,
       NOT_cpReq_363_BIT_36_924_932_AND_NOT_wci_busy__ETC___d3063,
       NOT_cpReq_363_BIT_36_924_932_AND_NOT_wci_busy__ETC___d3126,
       NOT_cpReq_363_BIT_36_924_932_AND_NOT_wci_busy__ETC___d3189,
       NOT_cpReq_363_BIT_36_924_932_AND_NOT_wci_busy__ETC___d3252,
       NOT_cpReq_363_BIT_36_924_932_AND_NOT_wci_busy__ETC___d3315,
       NOT_cpReq_363_BIT_36_924_932_AND_NOT_wci_busy__ETC___d3378,
       NOT_cpReq_363_BIT_36_924_932_AND_NOT_wci_busy__ETC___d3441,
       NOT_cpReq_363_BIT_36_924_932_AND_NOT_wci_busy__ETC___d3504,
       NOT_cpReq_363_BIT_36_924_932_AND_NOT_wci_busy__ETC___d3567,
       NOT_cpReq_363_BIT_36_924_932_AND_NOT_wci_busy__ETC___d3630,
       NOT_cpReq_363_BIT_36_924_932_AND_NOT_wci_busy__ETC___d3693,
       NOT_cpReq_363_BIT_36_924_932_AND_NOT_wci_busy__ETC___d3756,
       NOT_cpReq_363_BIT_36_924_932_AND_NOT_wci_busy__ETC___d3819,
       NOT_wci_busy_10_636_536_AND_wci_wReset_n_10_61_ETC___d3549,
       NOT_wci_busy_11_776_599_AND_wci_wReset_n_11_75_ETC___d3612,
       NOT_wci_busy_12_916_662_AND_wci_wReset_n_12_89_ETC___d3675,
       NOT_wci_busy_13_056_725_AND_wci_wReset_n_13_03_ETC___d3738,
       NOT_wci_busy_14_196_788_AND_wci_wReset_n_14_17_ETC___d3801,
       NOT_wci_busy_1_76_969_AND_wci_wReset_n_1_56_OR_ETC___d2982,
       NOT_wci_busy_2_16_032_AND_wci_wReset_n_2_96_OR_ETC___d3045,
       NOT_wci_busy_36_886_AND_wci_wReset_n_16_OR_wci_ETC___d2904,
       NOT_wci_busy_3_56_095_AND_wci_wReset_n_3_36_OR_ETC___d3108,
       NOT_wci_busy_4_96_158_AND_wci_wReset_n_4_76_OR_ETC___d3171,
       NOT_wci_busy_5_36_221_AND_wci_wReset_n_5_16_OR_ETC___d3234,
       NOT_wci_busy_6_076_284_AND_wci_wReset_n_6_056__ETC___d3297,
       NOT_wci_busy_7_216_347_AND_wci_wReset_n_7_196__ETC___d3360,
       NOT_wci_busy_8_356_410_AND_wci_wReset_n_8_336__ETC___d3423,
       NOT_wci_busy_9_496_473_AND_wci_wReset_n_9_476__ETC___d3486,
       cpReq_363_BITS_11_TO_4_366_EQ_0x30_595_OR_cpRe_ETC___d2632,
       cpReq_363_BITS_11_TO_4_366_ULT_0x30___d2438,
       cpReq_363_BITS_11_TO_4_366_ULT_0xC0___d2594,
       cpReq_363_BITS_27_TO_4_436_ULT_0x1000___d2866,
       cpReq_363_BITS_27_TO_4_436_ULT_0x100___d2437,
       cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_AND_NOT_w_ETC___d2953,
       cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_AND_NOT_w_ETC___d3019,
       cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_AND_NOT_w_ETC___d3082,
       cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_AND_NOT_w_ETC___d3145,
       cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_AND_NOT_w_ETC___d3208,
       cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_AND_NOT_w_ETC___d3271,
       cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_AND_NOT_w_ETC___d3334,
       cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_AND_NOT_w_ETC___d3397,
       cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_AND_NOT_w_ETC___d3460,
       cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_AND_NOT_w_ETC___d3523,
       cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_AND_NOT_w_ETC___d3586,
       cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_AND_NOT_w_ETC___d3649,
       cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_AND_NOT_w_ETC___d3712,
       cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_AND_NOT_w_ETC___d3775,
       cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_AND_NOT_w_ETC___d3838,
       cpReq_363_BIT_36_924_AND_NOT_wci_busy_10_636_5_ETC___d3560,
       cpReq_363_BIT_36_924_AND_NOT_wci_busy_11_776_5_ETC___d3623,
       cpReq_363_BIT_36_924_AND_NOT_wci_busy_12_916_6_ETC___d3686,
       cpReq_363_BIT_36_924_AND_NOT_wci_busy_13_056_7_ETC___d3749,
       cpReq_363_BIT_36_924_AND_NOT_wci_busy_14_196_7_ETC___d3812,
       cpReq_363_BIT_36_924_AND_NOT_wci_busy_1_76_969_ETC___d2993,
       cpReq_363_BIT_36_924_AND_NOT_wci_busy_2_16_032_ETC___d3056,
       cpReq_363_BIT_36_924_AND_NOT_wci_busy_36_886_A_ETC___d2925,
       cpReq_363_BIT_36_924_AND_NOT_wci_busy_3_56_095_ETC___d3119,
       cpReq_363_BIT_36_924_AND_NOT_wci_busy_4_96_158_ETC___d3182,
       cpReq_363_BIT_36_924_AND_NOT_wci_busy_5_36_221_ETC___d3245,
       cpReq_363_BIT_36_924_AND_NOT_wci_busy_6_076_28_ETC___d3308,
       cpReq_363_BIT_36_924_AND_NOT_wci_busy_7_216_34_ETC___d3371,
       cpReq_363_BIT_36_924_AND_NOT_wci_busy_8_356_41_ETC___d3434,
       cpReq_363_BIT_36_924_AND_NOT_wci_busy_9_496_47_ETC___d3497,
`ifdef not
       timeServ_ppsExtSync_d2_2_AND_NOT_timeServ_ppsE_ETC___d61,
       timeServ_ppsExtSync_d2_2_AND_NOT_timeServ_ppsE_ETC___d70,
       timeServ_refFromRise_3_ULE_199800000___d5459,
       timeServ_refFromRise_3_ULT_200200000___d5878,
`endif
       wci_respTimr_10_628_ULT_1_SL_wci_wTimeout_10_6_ETC___d5889,
       wci_respTimr_11_768_ULT_1_SL_wci_wTimeout_11_7_ETC___d5890,
       wci_respTimr_12_908_ULT_1_SL_wci_wTimeout_12_9_ETC___d5891,
       wci_respTimr_13_048_ULT_1_SL_wci_wTimeout_13_0_ETC___d5892,
       wci_respTimr_14_188_ULT_1_SL_wci_wTimeout_14_1_ETC___d5893,
       wci_respTimr_1_68_ULT_1_SL_wci_wTimeout_1_69_70___d5880,
       wci_respTimr_28_ULT_1_SL_wci_wTimeout_29_30___d5879,
       wci_respTimr_2_08_ULT_1_SL_wci_wTimeout_2_09_10___d5881,
       wci_respTimr_3_48_ULT_1_SL_wci_wTimeout_3_49_50___d5882,
       wci_respTimr_4_88_ULT_1_SL_wci_wTimeout_4_89_90___d5883,
       wci_respTimr_5_28_ULT_1_SL_wci_wTimeout_5_29_30___d5884,
       wci_respTimr_6_068_ULT_1_SL_wci_wTimeout_6_069_ETC___d5885,
       wci_respTimr_7_208_ULT_1_SL_wci_wTimeout_7_209_ETC___d5886,
       wci_respTimr_8_348_ULT_1_SL_wci_wTimeout_8_349_ETC___d5887,
       wci_respTimr_9_488_ULT_1_SL_wci_wTimeout_9_489_ETC___d5888,
       wci_wReset_n_10_616_AND_NOT_wci_busy_10_636_53_ETC___d3539,
       wci_wReset_n_11_756_AND_NOT_wci_busy_11_776_59_ETC___d3602,
       wci_wReset_n_12_896_AND_NOT_wci_busy_12_916_66_ETC___d3665,
       wci_wReset_n_13_036_AND_NOT_wci_busy_13_056_72_ETC___d3728,
       wci_wReset_n_14_176_AND_NOT_wci_busy_14_196_78_ETC___d3791,
       wci_wReset_n_16_AND_NOT_wci_busy_36_886_AND_NO_ETC___d2889,
       wci_wReset_n_1_56_AND_NOT_wci_busy_1_76_969_AN_ETC___d2972,
       wci_wReset_n_2_96_AND_NOT_wci_busy_2_16_032_AN_ETC___d3035,
       wci_wReset_n_3_36_AND_NOT_wci_busy_3_56_095_AN_ETC___d3098,
       wci_wReset_n_4_76_AND_NOT_wci_busy_4_96_158_AN_ETC___d3161,
       wci_wReset_n_5_16_AND_NOT_wci_busy_5_36_221_AN_ETC___d3224,
       wci_wReset_n_6_056_AND_NOT_wci_busy_6_076_284__ETC___d3287,
       wci_wReset_n_7_196_AND_NOT_wci_busy_7_216_347__ETC___d3350,
       wci_wReset_n_8_336_AND_NOT_wci_busy_8_356_410__ETC___d3413,
       wci_wReset_n_9_476_AND_NOT_wci_busy_9_496_473__ETC___d3476,
       wci_wciResponse_10_wget__623_BITS_33_TO_32_624_ETC___d1652,
       wci_wciResponse_11_wget__763_BITS_33_TO_32_764_ETC___d1792,
       wci_wciResponse_12_wget__903_BITS_33_TO_32_904_ETC___d1932,
       wci_wciResponse_13_wget__043_BITS_33_TO_32_044_ETC___d2072,
       wci_wciResponse_14_wget__183_BITS_33_TO_32_184_ETC___d2212,
       wci_wciResponse_1_wget__63_BITS_33_TO_32_64_EQ_ETC___d392,
       wci_wciResponse_2_wget__03_BITS_33_TO_32_04_EQ_ETC___d532,
       wci_wciResponse_3_wget__43_BITS_33_TO_32_44_EQ_ETC___d672,
       wci_wciResponse_4_wget__83_BITS_33_TO_32_84_EQ_ETC___d812,
       wci_wciResponse_5_wget__23_BITS_33_TO_32_24_EQ_ETC___d952,
       wci_wciResponse_6_wget__063_BITS_33_TO_32_064__ETC___d1092,
       wci_wciResponse_7_wget__203_BITS_33_TO_32_204__ETC___d1232,
       wci_wciResponse_8_wget__343_BITS_33_TO_32_344__ETC___d1372,
       wci_wciResponse_9_wget__483_BITS_33_TO_32_484__ETC___d1512,
       wci_wciResponse_wget__23_BITS_33_TO_32_24_EQ_0_ETC___d252;

  // output resets
  assign RST_N_wci_Vm_0 = wci_mReset$OUT_RST ;
  assign RST_N_wci_Vm_1 = wci_mReset_1$OUT_RST ;
  assign RST_N_wci_Vm_2 = wci_mReset_2$OUT_RST ;
  assign RST_N_wci_Vm_3 = wci_mReset_3$OUT_RST ;
  assign RST_N_wci_Vm_4 = wci_mReset_4$OUT_RST ;
  assign RST_N_wci_Vm_5 = wci_mReset_5$OUT_RST ;
  assign RST_N_wci_Vm_6 = wci_mReset_6$OUT_RST ;
  assign RST_N_wci_Vm_7 = wci_mReset_7$OUT_RST ;
  assign RST_N_wci_Vm_8 = wci_mReset_8$OUT_RST ;
  assign RST_N_wci_Vm_9 = wci_mReset_9$OUT_RST ;
  assign RST_N_wci_Vm_10 = wci_mReset_10$OUT_RST ;
  assign RST_N_wci_Vm_11 = wci_mReset_11$OUT_RST ;
  assign RST_N_wci_Vm_12 = wci_mReset_12$OUT_RST ;
  assign RST_N_wci_Vm_13 = wci_mReset_13$OUT_RST ;
  assign RST_N_wci_Vm_14 = wci_mReset_14$OUT_RST ;

  // action method server_request_put
  assign RDY_server_request_put = cpReqF$FULL_N ;

  // actionvalue method server_response_get
  assign server_response_get = cpRespF$D_OUT ;
  assign RDY_server_response_get = cpRespF$EMPTY_N ;

  // value method wci_Vm_0_mCmd
  assign wci_Vm_0_MCmd = wci_sThreadBusy_d ? 3'd0 : wci_reqF_q_0[71:69] ;

  // value method wci_Vm_0_mAddrSpace
  assign wci_Vm_0_MAddrSpace = !wci_sThreadBusy_d && wci_reqF_q_0[68] ;

  // value method wci_Vm_0_mByteEn
  assign wci_Vm_0_MByteEn = wci_sThreadBusy_d ? 4'd0 : wci_reqF_q_0[67:64] ;

  // value method wci_Vm_0_mAddr
  assign wci_Vm_0_MAddr = wci_sThreadBusy_d ? 32'd0 : wci_reqF_q_0[63:32] ;

  // value method wci_Vm_0_mData
  assign wci_Vm_0_MData = wci_reqF_q_0[31:0] ;

  // value method wci_Vm_0_mFlag
  assign wci_Vm_0_MFlag = wci_mFlagReg ;

  // value method wci_Vm_1_mCmd
  assign wci_Vm_1_MCmd = wci_sThreadBusy_d_1 ? 3'd0 : wci_reqF_1_q_0[71:69] ;

  // value method wci_Vm_1_mAddrSpace
  assign wci_Vm_1_MAddrSpace = !wci_sThreadBusy_d_1 && wci_reqF_1_q_0[68] ;

  // value method wci_Vm_1_mByteEn
  assign wci_Vm_1_MByteEn =
	     wci_sThreadBusy_d_1 ? 4'd0 : wci_reqF_1_q_0[67:64] ;

  // value method wci_Vm_1_mAddr
  assign wci_Vm_1_MAddr =
	     wci_sThreadBusy_d_1 ? 32'd0 : wci_reqF_1_q_0[63:32] ;

  // value method wci_Vm_1_mData
  assign wci_Vm_1_MData = wci_reqF_1_q_0[31:0] ;

  // value method wci_Vm_1_mFlag
  assign wci_Vm_1_MFlag = wci_mFlagReg_1 ;

  // value method wci_Vm_2_mCmd
  assign wci_Vm_2_MCmd = wci_sThreadBusy_d_2 ? 3'd0 : wci_reqF_2_q_0[71:69] ;

  // value method wci_Vm_2_mAddrSpace
  assign wci_Vm_2_MAddrSpace = !wci_sThreadBusy_d_2 && wci_reqF_2_q_0[68] ;

  // value method wci_Vm_2_mByteEn
  assign wci_Vm_2_MByteEn =
	     wci_sThreadBusy_d_2 ? 4'd0 : wci_reqF_2_q_0[67:64] ;

  // value method wci_Vm_2_mAddr
  assign wci_Vm_2_MAddr =
	     wci_sThreadBusy_d_2 ? 32'd0 : wci_reqF_2_q_0[63:32] ;

  // value method wci_Vm_2_mData
  assign wci_Vm_2_MData = wci_reqF_2_q_0[31:0] ;

  // value method wci_Vm_2_mFlag
  assign wci_Vm_2_MFlag = wci_mFlagReg_2 ;

  // value method wci_Vm_3_mCmd
  assign wci_Vm_3_MCmd = wci_sThreadBusy_d_3 ? 3'd0 : wci_reqF_3_q_0[71:69] ;

  // value method wci_Vm_3_mAddrSpace
  assign wci_Vm_3_MAddrSpace = !wci_sThreadBusy_d_3 && wci_reqF_3_q_0[68] ;

  // value method wci_Vm_3_mByteEn
  assign wci_Vm_3_MByteEn =
	     wci_sThreadBusy_d_3 ? 4'd0 : wci_reqF_3_q_0[67:64] ;

  // value method wci_Vm_3_mAddr
  assign wci_Vm_3_MAddr =
	     wci_sThreadBusy_d_3 ? 32'd0 : wci_reqF_3_q_0[63:32] ;

  // value method wci_Vm_3_mData
  assign wci_Vm_3_MData = wci_reqF_3_q_0[31:0] ;

  // value method wci_Vm_3_mFlag
  assign wci_Vm_3_MFlag = wci_mFlagReg_3 ;

  // value method wci_Vm_4_mCmd
  assign wci_Vm_4_MCmd = wci_sThreadBusy_d_4 ? 3'd0 : wci_reqF_4_q_0[71:69] ;

  // value method wci_Vm_4_mAddrSpace
  assign wci_Vm_4_MAddrSpace = !wci_sThreadBusy_d_4 && wci_reqF_4_q_0[68] ;

  // value method wci_Vm_4_mByteEn
  assign wci_Vm_4_MByteEn =
	     wci_sThreadBusy_d_4 ? 4'd0 : wci_reqF_4_q_0[67:64] ;

  // value method wci_Vm_4_mAddr
  assign wci_Vm_4_MAddr =
	     wci_sThreadBusy_d_4 ? 32'd0 : wci_reqF_4_q_0[63:32] ;

  // value method wci_Vm_4_mData
  assign wci_Vm_4_MData = wci_reqF_4_q_0[31:0] ;

  // value method wci_Vm_4_mFlag
  assign wci_Vm_4_MFlag = wci_mFlagReg_4 ;

  // value method wci_Vm_5_mCmd
  assign wci_Vm_5_MCmd = wci_sThreadBusy_d_5 ? 3'd0 : wci_reqF_5_q_0[71:69] ;

  // value method wci_Vm_5_mAddrSpace
  assign wci_Vm_5_MAddrSpace = !wci_sThreadBusy_d_5 && wci_reqF_5_q_0[68] ;

  // value method wci_Vm_5_mByteEn
  assign wci_Vm_5_MByteEn =
	     wci_sThreadBusy_d_5 ? 4'd0 : wci_reqF_5_q_0[67:64] ;

  // value method wci_Vm_5_mAddr
  assign wci_Vm_5_MAddr =
	     wci_sThreadBusy_d_5 ? 32'd0 : wci_reqF_5_q_0[63:32] ;

  // value method wci_Vm_5_mData
  assign wci_Vm_5_MData = wci_reqF_5_q_0[31:0] ;

  // value method wci_Vm_5_mFlag
  assign wci_Vm_5_MFlag = wci_mFlagReg_5 ;

  // value method wci_Vm_6_mCmd
  assign wci_Vm_6_MCmd = wci_sThreadBusy_d_6 ? 3'd0 : wci_reqF_6_q_0[71:69] ;

  // value method wci_Vm_6_mAddrSpace
  assign wci_Vm_6_MAddrSpace = !wci_sThreadBusy_d_6 && wci_reqF_6_q_0[68] ;

  // value method wci_Vm_6_mByteEn
  assign wci_Vm_6_MByteEn =
	     wci_sThreadBusy_d_6 ? 4'd0 : wci_reqF_6_q_0[67:64] ;

  // value method wci_Vm_6_mAddr
  assign wci_Vm_6_MAddr =
	     wci_sThreadBusy_d_6 ? 32'd0 : wci_reqF_6_q_0[63:32] ;

  // value method wci_Vm_6_mData
  assign wci_Vm_6_MData = wci_reqF_6_q_0[31:0] ;

  // value method wci_Vm_6_mFlag
  assign wci_Vm_6_MFlag = wci_mFlagReg_6 ;

  // value method wci_Vm_7_mCmd
  assign wci_Vm_7_MCmd = wci_sThreadBusy_d_7 ? 3'd0 : wci_reqF_7_q_0[71:69] ;

  // value method wci_Vm_7_mAddrSpace
  assign wci_Vm_7_MAddrSpace = !wci_sThreadBusy_d_7 && wci_reqF_7_q_0[68] ;

  // value method wci_Vm_7_mByteEn
  assign wci_Vm_7_MByteEn =
	     wci_sThreadBusy_d_7 ? 4'd0 : wci_reqF_7_q_0[67:64] ;

  // value method wci_Vm_7_mAddr
  assign wci_Vm_7_MAddr =
	     wci_sThreadBusy_d_7 ? 32'd0 : wci_reqF_7_q_0[63:32] ;

  // value method wci_Vm_7_mData
  assign wci_Vm_7_MData = wci_reqF_7_q_0[31:0] ;

  // value method wci_Vm_7_mFlag
  assign wci_Vm_7_MFlag = wci_mFlagReg_7 ;

  // value method wci_Vm_8_mCmd
  assign wci_Vm_8_MCmd = wci_sThreadBusy_d_8 ? 3'd0 : wci_reqF_8_q_0[71:69] ;

  // value method wci_Vm_8_mAddrSpace
  assign wci_Vm_8_MAddrSpace = !wci_sThreadBusy_d_8 && wci_reqF_8_q_0[68] ;

  // value method wci_Vm_8_mByteEn
  assign wci_Vm_8_MByteEn =
	     wci_sThreadBusy_d_8 ? 4'd0 : wci_reqF_8_q_0[67:64] ;

  // value method wci_Vm_8_mAddr
  assign wci_Vm_8_MAddr =
	     wci_sThreadBusy_d_8 ? 32'd0 : wci_reqF_8_q_0[63:32] ;

  // value method wci_Vm_8_mData
  assign wci_Vm_8_MData = wci_reqF_8_q_0[31:0] ;

  // value method wci_Vm_8_mFlag
  assign wci_Vm_8_MFlag = wci_mFlagReg_8 ;

  // value method wci_Vm_9_mCmd
  assign wci_Vm_9_MCmd = wci_sThreadBusy_d_9 ? 3'd0 : wci_reqF_9_q_0[71:69] ;

  // value method wci_Vm_9_mAddrSpace
  assign wci_Vm_9_MAddrSpace = !wci_sThreadBusy_d_9 && wci_reqF_9_q_0[68] ;

  // value method wci_Vm_9_mByteEn
  assign wci_Vm_9_MByteEn =
	     wci_sThreadBusy_d_9 ? 4'd0 : wci_reqF_9_q_0[67:64] ;

  // value method wci_Vm_9_mAddr
  assign wci_Vm_9_MAddr =
	     wci_sThreadBusy_d_9 ? 32'd0 : wci_reqF_9_q_0[63:32] ;

  // value method wci_Vm_9_mData
  assign wci_Vm_9_MData = wci_reqF_9_q_0[31:0] ;

  // value method wci_Vm_9_mFlag
  assign wci_Vm_9_MFlag = wci_mFlagReg_9 ;

  // value method wci_Vm_10_mCmd
  assign wci_Vm_10_MCmd =
	     wci_sThreadBusy_d_10 ? 3'd0 : wci_reqF_10_q_0[71:69] ;

  // value method wci_Vm_10_mAddrSpace
  assign wci_Vm_10_MAddrSpace = !wci_sThreadBusy_d_10 && wci_reqF_10_q_0[68] ;

  // value method wci_Vm_10_mByteEn
  assign wci_Vm_10_MByteEn =
	     wci_sThreadBusy_d_10 ? 4'd0 : wci_reqF_10_q_0[67:64] ;

  // value method wci_Vm_10_mAddr
  assign wci_Vm_10_MAddr =
	     wci_sThreadBusy_d_10 ? 32'd0 : wci_reqF_10_q_0[63:32] ;

  // value method wci_Vm_10_mData
  assign wci_Vm_10_MData = wci_reqF_10_q_0[31:0] ;

  // value method wci_Vm_10_mFlag
  assign wci_Vm_10_MFlag = wci_mFlagReg_10 ;

  // value method wci_Vm_11_mCmd
  assign wci_Vm_11_MCmd =
	     wci_sThreadBusy_d_11 ? 3'd0 : wci_reqF_11_q_0[71:69] ;

  // value method wci_Vm_11_mAddrSpace
  assign wci_Vm_11_MAddrSpace = !wci_sThreadBusy_d_11 && wci_reqF_11_q_0[68] ;

  // value method wci_Vm_11_mByteEn
  assign wci_Vm_11_MByteEn =
	     wci_sThreadBusy_d_11 ? 4'd0 : wci_reqF_11_q_0[67:64] ;

  // value method wci_Vm_11_mAddr
  assign wci_Vm_11_MAddr =
	     wci_sThreadBusy_d_11 ? 32'd0 : wci_reqF_11_q_0[63:32] ;

  // value method wci_Vm_11_mData
  assign wci_Vm_11_MData = wci_reqF_11_q_0[31:0] ;

  // value method wci_Vm_11_mFlag
  assign wci_Vm_11_MFlag = wci_mFlagReg_11 ;

  // value method wci_Vm_12_mCmd
  assign wci_Vm_12_MCmd =
	     wci_sThreadBusy_d_12 ? 3'd0 : wci_reqF_12_q_0[71:69] ;

  // value method wci_Vm_12_mAddrSpace
  assign wci_Vm_12_MAddrSpace = !wci_sThreadBusy_d_12 && wci_reqF_12_q_0[68] ;

  // value method wci_Vm_12_mByteEn
  assign wci_Vm_12_MByteEn =
	     wci_sThreadBusy_d_12 ? 4'd0 : wci_reqF_12_q_0[67:64] ;

  // value method wci_Vm_12_mAddr
  assign wci_Vm_12_MAddr =
	     wci_sThreadBusy_d_12 ? 32'd0 : wci_reqF_12_q_0[63:32] ;

  // value method wci_Vm_12_mData
  assign wci_Vm_12_MData = wci_reqF_12_q_0[31:0] ;

  // value method wci_Vm_12_mFlag
  assign wci_Vm_12_MFlag = wci_mFlagReg_12 ;

  // value method wci_Vm_13_mCmd
  assign wci_Vm_13_MCmd =
	     wci_sThreadBusy_d_13 ? 3'd0 : wci_reqF_13_q_0[71:69] ;

  // value method wci_Vm_13_mAddrSpace
  assign wci_Vm_13_MAddrSpace = !wci_sThreadBusy_d_13 && wci_reqF_13_q_0[68] ;

  // value method wci_Vm_13_mByteEn
  assign wci_Vm_13_MByteEn =
	     wci_sThreadBusy_d_13 ? 4'd0 : wci_reqF_13_q_0[67:64] ;

  // value method wci_Vm_13_mAddr
  assign wci_Vm_13_MAddr =
	     wci_sThreadBusy_d_13 ? 32'd0 : wci_reqF_13_q_0[63:32] ;

  // value method wci_Vm_13_mData
  assign wci_Vm_13_MData = wci_reqF_13_q_0[31:0] ;

  // value method wci_Vm_13_mFlag
  assign wci_Vm_13_MFlag = wci_mFlagReg_13 ;

  // value method wci_Vm_14_mCmd
  assign wci_Vm_14_MCmd =
	     wci_sThreadBusy_d_14 ? 3'd0 : wci_reqF_14_q_0[71:69] ;

  // value method wci_Vm_14_mAddrSpace
  assign wci_Vm_14_MAddrSpace = !wci_sThreadBusy_d_14 && wci_reqF_14_q_0[68] ;

  // value method wci_Vm_14_mByteEn
  assign wci_Vm_14_MByteEn =
	     wci_sThreadBusy_d_14 ? 4'd0 : wci_reqF_14_q_0[67:64] ;

  // value method wci_Vm_14_mAddr
  assign wci_Vm_14_MAddr =
	     wci_sThreadBusy_d_14 ? 32'd0 : wci_reqF_14_q_0[63:32] ;

  // value method wci_Vm_14_mData
  assign wci_Vm_14_MData = wci_reqF_14_q_0[31:0] ;

  // value method wci_Vm_14_mFlag
  assign wci_Vm_14_MFlag = wci_mFlagReg_14 ;

`ifdef not
  // value method cpNow
  assign cpNow = timeServ_now ;
  assign RDY_cpNow = 1'd1 ;

  // value method gps_ppsSyncOut
  always@(timeServ_ppsOutMode$dD_OUT or
	  timeServ_xo2 or timeServ_ppsDrive or timeServ_ppsExtSync_d2)
  begin
    case (timeServ_ppsOutMode$dD_OUT)
      2'd0: gps_ppsSyncOut = timeServ_ppsDrive;
      2'd1: gps_ppsSyncOut = timeServ_ppsExtSync_d2;
      default: gps_ppsSyncOut =
		   timeServ_ppsOutMode$dD_OUT == 2'd2 && timeServ_xo2;
    endcase
  end

  // value method led
  assign led = scratch24[1:0] ;
`endif

  // submodule adminResp1F
  FIFO1 #(.width(32'd33), .guarded(32'd1)) adminResp1F(.RST(RST_N),
						       .CLK(CLK),
						       .D_IN(adminResp1F$D_IN),
						       .ENQ(adminResp1F$ENQ),
						       .DEQ(adminResp1F$DEQ),
						       .CLR(adminResp1F$CLR),
						       .D_OUT(adminResp1F$D_OUT),
						       .FULL_N(adminResp1F$FULL_N),
						       .EMPTY_N(adminResp1F$EMPTY_N));

  // submodule adminResp2F
  FIFO1 #(.width(32'd33), .guarded(32'd1)) adminResp2F(.RST(RST_N),
						       .CLK(CLK),
						       .D_IN(adminResp2F$D_IN),
						       .ENQ(adminResp2F$ENQ),
						       .DEQ(adminResp2F$DEQ),
						       .CLR(adminResp2F$CLR),
						       .D_OUT(adminResp2F$D_OUT),
						       .FULL_N(adminResp2F$FULL_N),
						       .EMPTY_N(adminResp2F$EMPTY_N));

  // submodule adminResp3F
  FIFO1 #(.width(32'd33), .guarded(32'd1)) adminResp3F(.RST(RST_N),
						       .CLK(CLK),
						       .D_IN(adminResp3F$D_IN),
						       .ENQ(adminResp3F$ENQ),
						       .DEQ(adminResp3F$DEQ),
						       .CLR(adminResp3F$CLR),
						       .D_OUT(adminResp3F$D_OUT),
						       .FULL_N(adminResp3F$FULL_N),
						       .EMPTY_N(adminResp3F$EMPTY_N));

  // submodule adminResp4F
  FIFO1 #(.width(32'd33), .guarded(32'd1)) adminResp4F(.RST(RST_N),
						       .CLK(CLK),
						       .D_IN(adminResp4F$D_IN),
						       .ENQ(adminResp4F$ENQ),
						       .DEQ(adminResp4F$DEQ),
						       .CLR(adminResp4F$CLR),
						       .D_OUT(adminResp4F$D_OUT),
						       .FULL_N(adminResp4F$FULL_N),
						       .EMPTY_N(adminResp4F$EMPTY_N));

  // submodule adminRespF
  FIFO1 #(.width(32'd33), .guarded(32'd1)) adminRespF(.RST(RST_N),
						      .CLK(CLK),
						      .D_IN(adminRespF$D_IN),
						      .ENQ(adminRespF$ENQ),
						      .DEQ(adminRespF$DEQ),
						      .CLR(adminRespF$CLR),
						      .D_OUT(adminRespF$D_OUT),
						      .FULL_N(adminRespF$FULL_N),
						      .EMPTY_N(adminRespF$EMPTY_N));

  // submodule cpReqF
  FIFO2 #(.width(32'd59), .guarded(32'd1)) cpReqF(.RST(RST_N),
						  .CLK(CLK),
						  .D_IN(cpReqF$D_IN),
						  .ENQ(cpReqF$ENQ),
						  .DEQ(cpReqF$DEQ),
						  .CLR(cpReqF$CLR),
						  .D_OUT(cpReqF$D_OUT),
						  .FULL_N(cpReqF$FULL_N),
						  .EMPTY_N(cpReqF$EMPTY_N));

  // submodule cpRespF
  FIFO2 #(.width(32'd40), .guarded(32'd1)) cpRespF(.RST(RST_N),
						   .CLK(CLK),
						   .D_IN(cpRespF$D_IN),
						   .ENQ(cpRespF$ENQ),
						   .DEQ(cpRespF$DEQ),
						   .CLR(cpRespF$CLR),
						   .D_OUT(cpRespF$D_OUT),
						   .FULL_N(cpRespF$FULL_N),
						   .EMPTY_N(cpRespF$EMPTY_N));

`ifdef not
  // submodule dna_dna
  DNA_PORT dna_dna(.CLK(dna_dna$CLK),
		   .DIN(dna_dna$DIN),
		   .READ(dna_dna$READ),
		   .SHIFT(dna_dna$SHIFT),
		   .DOUT(dna_dna$DOUT));

  // submodule rom_serverAdapter_outDataCore
  SizedFIFO #(.p1width(32'd32),
	      .p2depth(32'd3),
	      .p3cntr_width(32'd1),
	      .guarded(32'd1)) rom_serverAdapter_outDataCore(.RST(RST_N),
							     .CLK(CLK),
							     .D_IN(rom_serverAdapter_outDataCore$D_IN),
							     .ENQ(rom_serverAdapter_outDataCore$ENQ),
							     .DEQ(rom_serverAdapter_outDataCore$DEQ),
							     .CLR(rom_serverAdapter_outDataCore$CLR),
							     .D_OUT(rom_serverAdapter_outDataCore$D_OUT),
							     .FULL_N(rom_serverAdapter_outDataCore$FULL_N),
							     .EMPTY_N(rom_serverAdapter_outDataCore$EMPTY_N));

  // submodule timeServ_disableServo
  SyncRegister #(.width(32'd1), .init(1'd0)) timeServ_disableServo(.sCLK(CLK),
								   .dCLK(CLK_time_clk),
								   .sRST(RST_N),
								   .sD_IN(timeServ_disableServo$sD_IN),
								   .sEN(timeServ_disableServo$sEN),
								   .dD_OUT(timeServ_disableServo$dD_OUT),
								   .sRDY(timeServ_disableServo$sRDY));

  // submodule timeServ_nowInCC
  SyncRegister #(.width(32'd64),
		 .init(64'd0)) timeServ_nowInCC(.sCLK(CLK_time_clk),
						.dCLK(CLK),
						.sRST(RST_N_time_rst),
						.sD_IN(timeServ_nowInCC$sD_IN),
						.sEN(timeServ_nowInCC$sEN),
						.dD_OUT(timeServ_nowInCC$dD_OUT),
						.sRDY(timeServ_nowInCC$sRDY));

  // submodule timeServ_ppsDisablePPS
  SyncRegister #(.width(32'd1),
		 .init(1'd0)) timeServ_ppsDisablePPS(.sCLK(CLK),
						     .dCLK(CLK_time_clk),
						     .sRST(RST_N),
						     .sD_IN(timeServ_ppsDisablePPS$sD_IN),
						     .sEN(timeServ_ppsDisablePPS$sEN),
						     .dD_OUT(timeServ_ppsDisablePPS$dD_OUT),
						     .sRDY(timeServ_ppsDisablePPS$sRDY));

  // submodule timeServ_ppsLostCC
  SyncRegister #(.width(32'd1),
		 .init(1'd0)) timeServ_ppsLostCC(.sCLK(CLK_time_clk),
						 .dCLK(CLK),
						 .sRST(RST_N_time_rst),
						 .sD_IN(timeServ_ppsLostCC$sD_IN),
						 .sEN(timeServ_ppsLostCC$sEN),
						 .dD_OUT(timeServ_ppsLostCC$dD_OUT),
						 .sRDY(timeServ_ppsLostCC$sRDY));

  // submodule timeServ_ppsOKCC
  SyncRegister #(.width(32'd1),
		 .init(1'd0)) timeServ_ppsOKCC(.sCLK(CLK_time_clk),
					       .dCLK(CLK),
					       .sRST(RST_N_time_rst),
					       .sD_IN(timeServ_ppsOKCC$sD_IN),
					       .sEN(timeServ_ppsOKCC$sEN),
					       .dD_OUT(timeServ_ppsOKCC$dD_OUT),
					       .sRDY(timeServ_ppsOKCC$sRDY));

  // submodule timeServ_ppsOutMode
  SyncRegister #(.width(32'd2), .init(2'd0)) timeServ_ppsOutMode(.sCLK(CLK),
								 .dCLK(CLK_time_clk),
								 .sRST(RST_N),
								 .sD_IN(timeServ_ppsOutMode$sD_IN),
								 .sEN(timeServ_ppsOutMode$sEN),
								 .dD_OUT(timeServ_ppsOutMode$dD_OUT),
								 .sRDY(timeServ_ppsOutMode$sRDY));

  // submodule timeServ_refPerPPS
  SyncRegister #(.width(32'd28),
		 .init(28'd0)) timeServ_refPerPPS(.sCLK(CLK_time_clk),
						  .dCLK(CLK),
						  .sRST(RST_N_time_rst),
						  .sD_IN(timeServ_refPerPPS$sD_IN),
						  .sEN(timeServ_refPerPPS$sEN),
						  .dD_OUT(timeServ_refPerPPS$dD_OUT),
						  .sRDY(timeServ_refPerPPS$sRDY));

  // submodule timeServ_rollingPPSIn
  SyncRegister #(.width(32'd8),
		 .init(8'd0)) timeServ_rollingPPSIn(.sCLK(CLK_time_clk),
						    .dCLK(CLK),
						    .sRST(RST_N_time_rst),
						    .sD_IN(timeServ_rollingPPSIn$sD_IN),
						    .sEN(timeServ_rollingPPSIn$sEN),
						    .dD_OUT(timeServ_rollingPPSIn$dD_OUT),
						    .sRDY(timeServ_rollingPPSIn$sRDY));

  // submodule timeServ_setRefF
  SyncFIFO #(.dataWidth(32'd64),
	     .depth(32'd2),
	     .indxWidth(32'd1)) timeServ_setRefF(.sCLK(CLK),
						 .dCLK(CLK_time_clk),
						 .sRST(RST_N),
						 .sD_IN(timeServ_setRefF$sD_IN),
						 .sENQ(timeServ_setRefF$sENQ),
						 .dDEQ(timeServ_setRefF$dDEQ),
						 .dD_OUT(timeServ_setRefF$dD_OUT),
						 .sFULL_N(timeServ_setRefF$sFULL_N),
						 .dEMPTY_N(timeServ_setRefF$dEMPTY_N));
`endif

  // submodule wci_mReset
  MakeResetA #(.RSTDELAY(32'd16), .init(1'd0)) wci_mReset(.CLK(CLK),
							  .RST(RST_N),
							  .DST_CLK(CLK),
							  .ASSERT_IN(wci_mReset$ASSERT_IN),
							  .ASSERT_OUT(),
							  .OUT_RST(wci_mReset$OUT_RST));

  // submodule wci_mReset_1
  MakeResetA #(.RSTDELAY(32'd16), .init(1'd0)) wci_mReset_1(.CLK(CLK),
							    .RST(RST_N),
							    .DST_CLK(CLK),
							    .ASSERT_IN(wci_mReset_1$ASSERT_IN),
							    .ASSERT_OUT(),
							    .OUT_RST(wci_mReset_1$OUT_RST));

  // submodule wci_mReset_10
  MakeResetA #(.RSTDELAY(32'd16), .init(1'd0)) wci_mReset_10(.CLK(CLK),
							     .RST(RST_N),
							     .DST_CLK(CLK),
							     .ASSERT_IN(wci_mReset_10$ASSERT_IN),
							     .ASSERT_OUT(),
							     .OUT_RST(wci_mReset_10$OUT_RST));

  // submodule wci_mReset_11
  MakeResetA #(.RSTDELAY(32'd16), .init(1'd0)) wci_mReset_11(.CLK(CLK),
							     .RST(RST_N),
							     .DST_CLK(CLK),
							     .ASSERT_IN(wci_mReset_11$ASSERT_IN),
							     .ASSERT_OUT(),
							     .OUT_RST(wci_mReset_11$OUT_RST));

  // submodule wci_mReset_12
  MakeResetA #(.RSTDELAY(32'd16), .init(1'd0)) wci_mReset_12(.CLK(CLK),
							     .RST(RST_N),
							     .DST_CLK(CLK),
							     .ASSERT_IN(wci_mReset_12$ASSERT_IN),
							     .ASSERT_OUT(),
							     .OUT_RST(wci_mReset_12$OUT_RST));

  // submodule wci_mReset_13
  MakeResetA #(.RSTDELAY(32'd16), .init(1'd0)) wci_mReset_13(.CLK(CLK),
							     .RST(RST_N),
							     .DST_CLK(CLK),
							     .ASSERT_IN(wci_mReset_13$ASSERT_IN),
							     .ASSERT_OUT(),
							     .OUT_RST(wci_mReset_13$OUT_RST));

  // submodule wci_mReset_14
  MakeResetA #(.RSTDELAY(32'd16), .init(1'd0)) wci_mReset_14(.CLK(CLK),
							     .RST(RST_N),
							     .DST_CLK(CLK),
							     .ASSERT_IN(wci_mReset_14$ASSERT_IN),
							     .ASSERT_OUT(),
							     .OUT_RST(wci_mReset_14$OUT_RST));

  // submodule wci_mReset_2
  MakeResetA #(.RSTDELAY(32'd16), .init(1'd0)) wci_mReset_2(.CLK(CLK),
							    .RST(RST_N),
							    .DST_CLK(CLK),
							    .ASSERT_IN(wci_mReset_2$ASSERT_IN),
							    .ASSERT_OUT(),
							    .OUT_RST(wci_mReset_2$OUT_RST));

  // submodule wci_mReset_3
  MakeResetA #(.RSTDELAY(32'd16), .init(1'd0)) wci_mReset_3(.CLK(CLK),
							    .RST(RST_N),
							    .DST_CLK(CLK),
							    .ASSERT_IN(wci_mReset_3$ASSERT_IN),
							    .ASSERT_OUT(),
							    .OUT_RST(wci_mReset_3$OUT_RST));

  // submodule wci_mReset_4
  MakeResetA #(.RSTDELAY(32'd16), .init(1'd0)) wci_mReset_4(.CLK(CLK),
							    .RST(RST_N),
							    .DST_CLK(CLK),
							    .ASSERT_IN(wci_mReset_4$ASSERT_IN),
							    .ASSERT_OUT(),
							    .OUT_RST(wci_mReset_4$OUT_RST));

  // submodule wci_mReset_5
  MakeResetA #(.RSTDELAY(32'd16), .init(1'd0)) wci_mReset_5(.CLK(CLK),
							    .RST(RST_N),
							    .DST_CLK(CLK),
							    .ASSERT_IN(wci_mReset_5$ASSERT_IN),
							    .ASSERT_OUT(),
							    .OUT_RST(wci_mReset_5$OUT_RST));

  // submodule wci_mReset_6
  MakeResetA #(.RSTDELAY(32'd16), .init(1'd0)) wci_mReset_6(.CLK(CLK),
							    .RST(RST_N),
							    .DST_CLK(CLK),
							    .ASSERT_IN(wci_mReset_6$ASSERT_IN),
							    .ASSERT_OUT(),
							    .OUT_RST(wci_mReset_6$OUT_RST));

  // submodule wci_mReset_7
  MakeResetA #(.RSTDELAY(32'd16), .init(1'd0)) wci_mReset_7(.CLK(CLK),
							    .RST(RST_N),
							    .DST_CLK(CLK),
							    .ASSERT_IN(wci_mReset_7$ASSERT_IN),
							    .ASSERT_OUT(),
							    .OUT_RST(wci_mReset_7$OUT_RST));

  // submodule wci_mReset_8
  MakeResetA #(.RSTDELAY(32'd16), .init(1'd0)) wci_mReset_8(.CLK(CLK),
							    .RST(RST_N),
							    .DST_CLK(CLK),
							    .ASSERT_IN(wci_mReset_8$ASSERT_IN),
							    .ASSERT_OUT(),
							    .OUT_RST(wci_mReset_8$OUT_RST));

  // submodule wci_mReset_9
  MakeResetA #(.RSTDELAY(32'd16), .init(1'd0)) wci_mReset_9(.CLK(CLK),
							    .RST(RST_N),
							    .DST_CLK(CLK),
							    .ASSERT_IN(wci_mReset_9$ASSERT_IN),
							    .ASSERT_OUT(),
							    .OUT_RST(wci_mReset_9$OUT_RST));

  // submodule wci_respF
  FIFO1 #(.width(32'd34), .guarded(32'd1)) wci_respF(.RST(RST_N),
						     .CLK(CLK),
						     .D_IN(wci_respF$D_IN),
						     .ENQ(wci_respF$ENQ),
						     .DEQ(wci_respF$DEQ),
						     .CLR(wci_respF$CLR),
						     .D_OUT(wci_respF$D_OUT),
						     .FULL_N(wci_respF$FULL_N),
						     .EMPTY_N(wci_respF$EMPTY_N));

  // submodule wci_respF_1
  FIFO1 #(.width(32'd34), .guarded(32'd1)) wci_respF_1(.RST(RST_N),
						       .CLK(CLK),
						       .D_IN(wci_respF_1$D_IN),
						       .ENQ(wci_respF_1$ENQ),
						       .DEQ(wci_respF_1$DEQ),
						       .CLR(wci_respF_1$CLR),
						       .D_OUT(wci_respF_1$D_OUT),
						       .FULL_N(wci_respF_1$FULL_N),
						       .EMPTY_N(wci_respF_1$EMPTY_N));

  // submodule wci_respF_10
  FIFO1 #(.width(32'd34), .guarded(32'd1)) wci_respF_10(.RST(RST_N),
							.CLK(CLK),
							.D_IN(wci_respF_10$D_IN),
							.ENQ(wci_respF_10$ENQ),
							.DEQ(wci_respF_10$DEQ),
							.CLR(wci_respF_10$CLR),
							.D_OUT(wci_respF_10$D_OUT),
							.FULL_N(wci_respF_10$FULL_N),
							.EMPTY_N(wci_respF_10$EMPTY_N));

  // submodule wci_respF_11
  FIFO1 #(.width(32'd34), .guarded(32'd1)) wci_respF_11(.RST(RST_N),
							.CLK(CLK),
							.D_IN(wci_respF_11$D_IN),
							.ENQ(wci_respF_11$ENQ),
							.DEQ(wci_respF_11$DEQ),
							.CLR(wci_respF_11$CLR),
							.D_OUT(wci_respF_11$D_OUT),
							.FULL_N(wci_respF_11$FULL_N),
							.EMPTY_N(wci_respF_11$EMPTY_N));

  // submodule wci_respF_12
  FIFO1 #(.width(32'd34), .guarded(32'd1)) wci_respF_12(.RST(RST_N),
							.CLK(CLK),
							.D_IN(wci_respF_12$D_IN),
							.ENQ(wci_respF_12$ENQ),
							.DEQ(wci_respF_12$DEQ),
							.CLR(wci_respF_12$CLR),
							.D_OUT(wci_respF_12$D_OUT),
							.FULL_N(wci_respF_12$FULL_N),
							.EMPTY_N(wci_respF_12$EMPTY_N));

  // submodule wci_respF_13
  FIFO1 #(.width(32'd34), .guarded(32'd1)) wci_respF_13(.RST(RST_N),
							.CLK(CLK),
							.D_IN(wci_respF_13$D_IN),
							.ENQ(wci_respF_13$ENQ),
							.DEQ(wci_respF_13$DEQ),
							.CLR(wci_respF_13$CLR),
							.D_OUT(wci_respF_13$D_OUT),
							.FULL_N(wci_respF_13$FULL_N),
							.EMPTY_N(wci_respF_13$EMPTY_N));

  // submodule wci_respF_14
  FIFO1 #(.width(32'd34), .guarded(32'd1)) wci_respF_14(.RST(RST_N),
							.CLK(CLK),
							.D_IN(wci_respF_14$D_IN),
							.ENQ(wci_respF_14$ENQ),
							.DEQ(wci_respF_14$DEQ),
							.CLR(wci_respF_14$CLR),
							.D_OUT(wci_respF_14$D_OUT),
							.FULL_N(wci_respF_14$FULL_N),
							.EMPTY_N(wci_respF_14$EMPTY_N));

  // submodule wci_respF_2
  FIFO1 #(.width(32'd34), .guarded(32'd1)) wci_respF_2(.RST(RST_N),
						       .CLK(CLK),
						       .D_IN(wci_respF_2$D_IN),
						       .ENQ(wci_respF_2$ENQ),
						       .DEQ(wci_respF_2$DEQ),
						       .CLR(wci_respF_2$CLR),
						       .D_OUT(wci_respF_2$D_OUT),
						       .FULL_N(wci_respF_2$FULL_N),
						       .EMPTY_N(wci_respF_2$EMPTY_N));

  // submodule wci_respF_3
  FIFO1 #(.width(32'd34), .guarded(32'd1)) wci_respF_3(.RST(RST_N),
						       .CLK(CLK),
						       .D_IN(wci_respF_3$D_IN),
						       .ENQ(wci_respF_3$ENQ),
						       .DEQ(wci_respF_3$DEQ),
						       .CLR(wci_respF_3$CLR),
						       .D_OUT(wci_respF_3$D_OUT),
						       .FULL_N(wci_respF_3$FULL_N),
						       .EMPTY_N(wci_respF_3$EMPTY_N));

  // submodule wci_respF_4
  FIFO1 #(.width(32'd34), .guarded(32'd1)) wci_respF_4(.RST(RST_N),
						       .CLK(CLK),
						       .D_IN(wci_respF_4$D_IN),
						       .ENQ(wci_respF_4$ENQ),
						       .DEQ(wci_respF_4$DEQ),
						       .CLR(wci_respF_4$CLR),
						       .D_OUT(wci_respF_4$D_OUT),
						       .FULL_N(wci_respF_4$FULL_N),
						       .EMPTY_N(wci_respF_4$EMPTY_N));

  // submodule wci_respF_5
  FIFO1 #(.width(32'd34), .guarded(32'd1)) wci_respF_5(.RST(RST_N),
						       .CLK(CLK),
						       .D_IN(wci_respF_5$D_IN),
						       .ENQ(wci_respF_5$ENQ),
						       .DEQ(wci_respF_5$DEQ),
						       .CLR(wci_respF_5$CLR),
						       .D_OUT(wci_respF_5$D_OUT),
						       .FULL_N(wci_respF_5$FULL_N),
						       .EMPTY_N(wci_respF_5$EMPTY_N));

  // submodule wci_respF_6
  FIFO1 #(.width(32'd34), .guarded(32'd1)) wci_respF_6(.RST(RST_N),
						       .CLK(CLK),
						       .D_IN(wci_respF_6$D_IN),
						       .ENQ(wci_respF_6$ENQ),
						       .DEQ(wci_respF_6$DEQ),
						       .CLR(wci_respF_6$CLR),
						       .D_OUT(wci_respF_6$D_OUT),
						       .FULL_N(wci_respF_6$FULL_N),
						       .EMPTY_N(wci_respF_6$EMPTY_N));

  // submodule wci_respF_7
  FIFO1 #(.width(32'd34), .guarded(32'd1)) wci_respF_7(.RST(RST_N),
						       .CLK(CLK),
						       .D_IN(wci_respF_7$D_IN),
						       .ENQ(wci_respF_7$ENQ),
						       .DEQ(wci_respF_7$DEQ),
						       .CLR(wci_respF_7$CLR),
						       .D_OUT(wci_respF_7$D_OUT),
						       .FULL_N(wci_respF_7$FULL_N),
						       .EMPTY_N(wci_respF_7$EMPTY_N));

  // submodule wci_respF_8
  FIFO1 #(.width(32'd34), .guarded(32'd1)) wci_respF_8(.RST(RST_N),
						       .CLK(CLK),
						       .D_IN(wci_respF_8$D_IN),
						       .ENQ(wci_respF_8$ENQ),
						       .DEQ(wci_respF_8$DEQ),
						       .CLR(wci_respF_8$CLR),
						       .D_OUT(wci_respF_8$D_OUT),
						       .FULL_N(wci_respF_8$FULL_N),
						       .EMPTY_N(wci_respF_8$EMPTY_N));

  // submodule wci_respF_9
  FIFO1 #(.width(32'd34), .guarded(32'd1)) wci_respF_9(.RST(RST_N),
						       .CLK(CLK),
						       .D_IN(wci_respF_9$D_IN),
						       .ENQ(wci_respF_9$ENQ),
						       .DEQ(wci_respF_9$DEQ),
						       .CLR(wci_respF_9$CLR),
						       .D_OUT(wci_respF_9$D_OUT),
						       .FULL_N(wci_respF_9$FULL_N),
						       .EMPTY_N(wci_respF_9$EMPTY_N));

  // rule RL_readAdminResponseCollect
  assign WILL_FIRE_RL_readAdminResponseCollect =
	     adminResp1F$EMPTY_N ?
	       adminRespF$FULL_N && adminResp1F$EMPTY_N :
	       (adminResp2F$EMPTY_N ?
		  adminRespF$FULL_N && adminResp2F$EMPTY_N :
		  (adminResp3F$EMPTY_N ?
		     adminRespF$FULL_N && adminResp3F$EMPTY_N :
		     !adminResp4F$EMPTY_N || adminRespF$FULL_N)) ;

  // rule RL_cpDispatch_T_T
  assign WILL_FIRE_RL_cpDispatch_T_T =
	     cpReq[64:62] == 3'd1 && cpReq[11:4] == 8'h20 && !dispatched ;

  // rule RL_cpDispatch_T_F_T
  assign WILL_FIRE_RL_cpDispatch_T_F_T =
	     cpReq[64:62] == 3'd1 && cpReq[11:4] == 8'h24 && !dispatched ;

  // rule RL_cpDispatch_T_F_F_T
  assign WILL_FIRE_RL_cpDispatch_T_F_F_T =
	     cpReq[64:62] == 3'd1 && cpReq[11:4] == 8'h28 && !dispatched ;

  // rule RL_cpDispatch_T_F_F_F_T
  assign WILL_FIRE_RL_cpDispatch_T_F_F_F_T =
	     cpReq[64:62] == 3'd1 && cpReq[11:4] == 8'h2C && !dispatched ;

  // rule RL_cpDispatch_T_F_F_F_F_F_T
  assign WILL_FIRE_RL_cpDispatch_T_F_F_F_F_F_T =
	     cpReq[64:62] == 3'd1 && cpReq[11:4] == 8'h38 && !dispatched ;

  // rule RL_cpDispatch_T_F_F_F_F_F_F_T
  assign WILL_FIRE_RL_cpDispatch_T_F_F_F_F_F_F_T =
`ifdef not
	     cpReq[64:62] == 3'd1 && cpReq[11:4] == 8'h3C &&
	     timeServ_setRefF$sFULL_N &&
	     !dispatched ;
`else
	      0;
`endif
  // rule RL_cpDispatch_T_F_F_F_F_F_F_F_T
  assign WILL_FIRE_RL_cpDispatch_T_F_F_F_F_F_F_F_T =
	     cpReq[64:62] == 3'd1 && cpReq[11:4] == 8'h40 && !dispatched ;

  // rule RL_cpDispatch_T_F_F_F_F_F_F_F_F_T
  assign WILL_FIRE_RL_cpDispatch_T_F_F_F_F_F_F_F_F_T =
	     cpReq[64:62] == 3'd1 && cpReq[11:4] == 8'h44 && !dispatched ;

  // rule RL_cpDispatch_T_F_F_F_F_F_F_F_F_F_T
  assign WILL_FIRE_RL_cpDispatch_T_F_F_F_F_F_F_F_F_F_T =
	     cpReq[64:62] == 3'd1 && cpReq[11:4] == 8'h4C && !dispatched ;

  // rule RL_cpDispatch_T_F_F_F_F_F_F_F_F_F_F
  assign WILL_FIRE_RL_cpDispatch_T_F_F_F_F_F_F_F_F_F_F =
	     cpReq[64:62] == 3'd1 && cpReq[11:4] != 8'h20 &&
	     cpReq[11:4] != 8'h24 &&
	     cpReq[11:4] != 8'h28 &&
	     cpReq[11:4] != 8'h2C &&
	     cpReq[11:4] != 8'h34 &&
	     cpReq[11:4] != 8'h38 &&
	     cpReq[11:4] != 8'h3C &&
	     cpReq[11:4] != 8'h40 &&
	     cpReq[11:4] != 8'h44 &&
	     cpReq[11:4] != 8'h4C &&
	     !dispatched ;

  // rule RL_cpDispatch_F_T_T_T
  assign CAN_FIRE_RL_cpDispatch_F_T_T_T =
	     cpReq[64:62] == 3'd2 &&
	     cpReq_363_BITS_27_TO_4_436_ULT_0x100___d2437 &&
	     cpReq_363_BITS_11_TO_4_366_ULT_0x30___d2438 &&
	     adminResp1F$FULL_N &&
	     !dispatched ;
  assign WILL_FIRE_RL_cpDispatch_F_T_T_T =
	     CAN_FIRE_RL_cpDispatch_F_T_T_T && !WILL_FIRE_RL_responseAdminRd ;

  // rule RL_cpDispatch_F_T_T_F_T_T
  assign CAN_FIRE_RL_cpDispatch_F_T_T_F_T_T =
	     cpReq[64:62] == 3'd2 &&
	     cpReq_363_BITS_27_TO_4_436_ULT_0x100___d2437 &&
	     !cpReq_363_BITS_11_TO_4_366_ULT_0x30___d2438 &&
	     cpReq_363_BITS_11_TO_4_366_ULT_0xC0___d2594 &&
	     cpReq_363_BITS_11_TO_4_366_EQ_0x30_595_OR_cpRe_ETC___d2632 ;
  assign WILL_FIRE_RL_cpDispatch_F_T_T_F_T_T =
	     CAN_FIRE_RL_cpDispatch_F_T_T_F_T_T &&
	     !WILL_FIRE_RL_responseAdminRd ;

  // rule RL_cpDispatch_F_T_T_F_T_F_T
  assign CAN_FIRE_RL_cpDispatch_F_T_T_F_T_F_T =
	     cpReq[64:62] == 3'd2 &&
	     cpReq_363_BITS_27_TO_4_436_ULT_0x100___d2437 &&
	     !cpReq_363_BITS_11_TO_4_366_ULT_0x30___d2438 &&
	     cpReq_363_BITS_11_TO_4_366_ULT_0xC0___d2594 &&
	     cpReq[11:4] == 8'h4C &&
	     adminResp2F$FULL_N &&
	     !dispatched ;
  assign WILL_FIRE_RL_cpDispatch_F_T_T_F_T_F_T =
	     CAN_FIRE_RL_cpDispatch_F_T_T_F_T_F_T &&
	     !WILL_FIRE_RL_responseAdminRd ;

  // rule RL_cpDispatch_F_T_T_F_T_F_F
  assign CAN_FIRE_RL_cpDispatch_F_T_T_F_T_F_F =
	     cpReq[64:62] == 3'd2 &&
	     cpReq_363_BITS_27_TO_4_436_ULT_0x100___d2437 &&
	     !cpReq_363_BITS_11_TO_4_366_ULT_0x30___d2438 &&
	     cpReq_363_BITS_11_TO_4_366_ULT_0xC0___d2594 &&
	     NOT_cpReq_363_BITS_11_TO_4_366_EQ_0x30_595_649_ETC___d2712 ;
  assign WILL_FIRE_RL_cpDispatch_F_T_T_F_T_F_F =
	     CAN_FIRE_RL_cpDispatch_F_T_T_F_T_F_F &&
	     !WILL_FIRE_RL_responseAdminRd ;

  // rule RL_cpDispatch_F_T_T_F_F
  assign CAN_FIRE_RL_cpDispatch_F_T_T_F_F =
	     cpReq[64:62] == 3'd2 &&
	     cpReq_363_BITS_27_TO_4_436_ULT_0x100___d2437 &&
	     !cpReq_363_BITS_11_TO_4_366_ULT_0x30___d2438 &&
	     !cpReq_363_BITS_11_TO_4_366_ULT_0xC0___d2594 &&
	     adminResp3F$FULL_N &&
	     !dispatched ;
  assign WILL_FIRE_RL_cpDispatch_F_T_T_F_F =
	     CAN_FIRE_RL_cpDispatch_F_T_T_F_F &&
	     !WILL_FIRE_RL_responseAdminRd ;

  // rule RL_cpDispatch_F_T_F_T
  assign WILL_FIRE_RL_cpDispatch_F_T_F_T =
	     cpReq[64:62] == 3'd2 &&
	     !cpReq_363_BITS_27_TO_4_436_ULT_0x100___d2437 &&
	     cpReq_363_BITS_27_TO_4_436_ULT_0x1000___d2866 &&
	     !dispatched &&
	     !WILL_FIRE_RL_responseAdminRd ;

`ifdef not
  // rule RL_cpDispatch_F_T_F_F
  assign CAN_FIRE_RL_cpDispatch_F_T_F_F =
	     cpReq[64:62] == 3'd2 &&
	     !cpReq_363_BITS_27_TO_4_436_ULT_0x100___d2437 &&
	     !cpReq_363_BITS_27_TO_4_436_ULT_0x1000___d2866 &&
	     (rom_serverAdapter_cnt ^ 3'h4) < 3'd7 &&
	     !dispatched ;
`endif
  // rule RL_cpDispatch_F_F_T_T_T_F
  assign WILL_FIRE_RL_cpDispatch_F_F_T_T_T_F =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd0 &&
	     cpReq[61:60] == 2'd2 &&
	     !wci_wReset_n &&
	     NOT_wci_busy_36_886_AND_wci_wReset_n_16_OR_wci_ETC___d2904 ;

  // rule RL_cpDispatch_F_F_T_T_F_T
  assign WILL_FIRE_RL_cpDispatch_F_F_T_T_F_T =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd0 &&
	     cpReq[61:60] == 2'd1 &&
	     cpReq[19:9] == 11'd0 &&
	     !wci_busy &&
	     wci_respF$FULL_N &&
	     !dispatched ;

  // rule RL_cpDispatch_F_F_T_T_F_F_F_T
  assign WILL_FIRE_RL_cpDispatch_F_F_T_T_F_F_F_T =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd0 &&
	     cpReq[61:60] != 2'd2 &&
	     (cpReq[61:60] != 2'd1 || cpReq[19:9] != 11'd0) &&
	     cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_AND_NOT_w_ETC___d2953 ;

  // rule RL_cpDispatch_F_F_T_T_F_F_F_F
  assign WILL_FIRE_RL_cpDispatch_F_F_T_T_F_F_F_F =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd0 &&
	     cpReq[61:60] != 2'd2 &&
	     (cpReq[61:60] != 2'd1 || cpReq[19:9] != 11'd0) &&
	     cpReq[9:6] != 4'h9 &&
	     NOT_cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_961_A_ETC___d2962 ;

  // rule RL_cpDispatch_F_F_T_F_T_T_F
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_T_T_F =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd1 &&
	     cpReq[61:60] == 2'd2 &&
	     !wci_wReset_n_1 &&
	     NOT_wci_busy_1_76_969_AND_wci_wReset_n_1_56_OR_ETC___d2982 ;

  // rule RL_cpDispatch_F_F_T_F_T_F_T
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_T_F_T =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd1 &&
	     cpReq[61:60] == 2'd1 &&
	     cpReq[19:9] == 11'd0 &&
	     !wci_busy_1 &&
	     wci_respF_1$FULL_N &&
	     !dispatched ;

  // rule RL_cpDispatch_F_F_T_F_T_F_F_F_T
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_T_F_F_F_T =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd1 &&
	     cpReq[61:60] != 2'd2 &&
	     (cpReq[61:60] != 2'd1 || cpReq[19:9] != 11'd0) &&
	     cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_AND_NOT_w_ETC___d3019 ;

  // rule RL_cpDispatch_F_F_T_F_T_F_F_F_F
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_T_F_F_F_F =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd1 &&
	     cpReq[61:60] != 2'd2 &&
	     (cpReq[61:60] != 2'd1 || cpReq[19:9] != 11'd0) &&
	     cpReq[9:6] != 4'h9 &&
	     NOT_cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_961_A_ETC___d3025 ;

  // rule RL_cpDispatch_F_F_T_F_F_T_T_F
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_T_F =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd2 &&
	     cpReq[61:60] == 2'd2 &&
	     !wci_wReset_n_2 &&
	     NOT_wci_busy_2_16_032_AND_wci_wReset_n_2_96_OR_ETC___d3045 ;

  // rule RL_cpDispatch_F_F_T_F_F_T_F_T
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_F_T =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd2 &&
	     cpReq[61:60] == 2'd1 &&
	     cpReq[19:9] == 11'd0 &&
	     !wci_busy_2 &&
	     wci_respF_2$FULL_N &&
	     !dispatched ;

  // rule RL_cpDispatch_F_F_T_F_F_T_F_F_F_T
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_F_F_F_T =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd2 &&
	     cpReq[61:60] != 2'd2 &&
	     (cpReq[61:60] != 2'd1 || cpReq[19:9] != 11'd0) &&
	     cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_AND_NOT_w_ETC___d3082 ;

  // rule RL_cpDispatch_F_F_T_F_F_T_F_F_F_F
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_F_F_F_F =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd2 &&
	     cpReq[61:60] != 2'd2 &&
	     (cpReq[61:60] != 2'd1 || cpReq[19:9] != 11'd0) &&
	     cpReq[9:6] != 4'h9 &&
	     NOT_cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_961_A_ETC___d3088 ;

  // rule RL_cpDispatch_F_F_T_F_F_F_T_T_F
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_T_F =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd3 &&
	     cpReq[61:60] == 2'd2 &&
	     !wci_wReset_n_3 &&
	     NOT_wci_busy_3_56_095_AND_wci_wReset_n_3_36_OR_ETC___d3108 ;

  // rule RL_cpDispatch_F_F_T_F_F_F_T_F_T
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_F_T =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd3 &&
	     cpReq[61:60] == 2'd1 &&
	     cpReq[19:9] == 11'd0 &&
	     !wci_busy_3 &&
	     wci_respF_3$FULL_N &&
	     !dispatched ;

  // rule RL_cpDispatch_F_F_T_F_F_F_T_F_F_F_T
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_F_F_F_T =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd3 &&
	     cpReq[61:60] != 2'd2 &&
	     (cpReq[61:60] != 2'd1 || cpReq[19:9] != 11'd0) &&
	     cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_AND_NOT_w_ETC___d3145 ;

  // rule RL_cpDispatch_F_F_T_F_F_F_T_F_F_F_F
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_F_F_F_F =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd3 &&
	     cpReq[61:60] != 2'd2 &&
	     (cpReq[61:60] != 2'd1 || cpReq[19:9] != 11'd0) &&
	     cpReq[9:6] != 4'h9 &&
	     NOT_cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_961_A_ETC___d3151 ;

  // rule RL_cpDispatch_F_F_T_F_F_F_F_T_T_F
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_T_F =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd4 &&
	     cpReq[61:60] == 2'd2 &&
	     !wci_wReset_n_4 &&
	     NOT_wci_busy_4_96_158_AND_wci_wReset_n_4_76_OR_ETC___d3171 ;

  // rule RL_cpDispatch_F_F_T_F_F_F_F_T_F_T
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_F_T =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd4 &&
	     cpReq[61:60] == 2'd1 &&
	     cpReq[19:9] == 11'd0 &&
	     !wci_busy_4 &&
	     wci_respF_4$FULL_N &&
	     !dispatched ;

  // rule RL_cpDispatch_F_F_T_F_F_F_F_T_F_F_F_T
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_F_F_F_T =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd4 &&
	     cpReq[61:60] != 2'd2 &&
	     (cpReq[61:60] != 2'd1 || cpReq[19:9] != 11'd0) &&
	     cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_AND_NOT_w_ETC___d3208 ;

  // rule RL_cpDispatch_F_F_T_F_F_F_F_T_F_F_F_F
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_F_F_F_F =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd4 &&
	     cpReq[61:60] != 2'd2 &&
	     (cpReq[61:60] != 2'd1 || cpReq[19:9] != 11'd0) &&
	     cpReq[9:6] != 4'h9 &&
	     NOT_cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_961_A_ETC___d3214 ;

  // rule RL_cpDispatch_F_F_T_F_F_F_F_F_T_T_F
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_T_F =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd5 &&
	     cpReq[61:60] == 2'd2 &&
	     !wci_wReset_n_5 &&
	     NOT_wci_busy_5_36_221_AND_wci_wReset_n_5_16_OR_ETC___d3234 ;

  // rule RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_T
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_T =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd5 &&
	     cpReq[61:60] == 2'd1 &&
	     cpReq[19:9] == 11'd0 &&
	     !wci_busy_5 &&
	     wci_respF_5$FULL_N &&
	     !dispatched ;

  // rule RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_F_F_T
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_F_F_T =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd5 &&
	     cpReq[61:60] != 2'd2 &&
	     (cpReq[61:60] != 2'd1 || cpReq[19:9] != 11'd0) &&
	     cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_AND_NOT_w_ETC___d3271 ;

  // rule RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_F_F_F
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_F_F_F =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd5 &&
	     cpReq[61:60] != 2'd2 &&
	     (cpReq[61:60] != 2'd1 || cpReq[19:9] != 11'd0) &&
	     cpReq[9:6] != 4'h9 &&
	     NOT_cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_961_A_ETC___d3277 ;

  // rule RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_T_F
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_T_F =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd6 &&
	     cpReq[61:60] == 2'd2 &&
	     !wci_wReset_n_6 &&
	     NOT_wci_busy_6_076_284_AND_wci_wReset_n_6_056__ETC___d3297 ;

  // rule RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_T
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_T =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd6 &&
	     cpReq[61:60] == 2'd1 &&
	     cpReq[19:9] == 11'd0 &&
	     !wci_busy_6 &&
	     wci_respF_6$FULL_N &&
	     !dispatched ;

  // rule RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_F_F_T
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_F_F_T =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd6 &&
	     cpReq[61:60] != 2'd2 &&
	     (cpReq[61:60] != 2'd1 || cpReq[19:9] != 11'd0) &&
	     cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_AND_NOT_w_ETC___d3334 ;

  // rule RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_F_F_F
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_F_F_F =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd6 &&
	     cpReq[61:60] != 2'd2 &&
	     (cpReq[61:60] != 2'd1 || cpReq[19:9] != 11'd0) &&
	     cpReq[9:6] != 4'h9 &&
	     NOT_cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_961_A_ETC___d3340 ;

  // rule RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_T_F
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_T_F =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd7 &&
	     cpReq[61:60] == 2'd2 &&
	     !wci_wReset_n_7 &&
	     NOT_wci_busy_7_216_347_AND_wci_wReset_n_7_196__ETC___d3360 ;

  // rule RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_T
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_T =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd7 &&
	     cpReq[61:60] == 2'd1 &&
	     cpReq[19:9] == 11'd0 &&
	     !wci_busy_7 &&
	     wci_respF_7$FULL_N &&
	     !dispatched ;

  // rule RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_F_F_T
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_F_F_T =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd7 &&
	     cpReq[61:60] != 2'd2 &&
	     (cpReq[61:60] != 2'd1 || cpReq[19:9] != 11'd0) &&
	     cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_AND_NOT_w_ETC___d3397 ;

  // rule RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_F_F_F
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_F_F_F =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd7 &&
	     cpReq[61:60] != 2'd2 &&
	     (cpReq[61:60] != 2'd1 || cpReq[19:9] != 11'd0) &&
	     cpReq[9:6] != 4'h9 &&
	     NOT_cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_961_A_ETC___d3403 ;

  // rule RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_T_F
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_T_F =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd8 &&
	     cpReq[61:60] == 2'd2 &&
	     !wci_wReset_n_8 &&
	     NOT_wci_busy_8_356_410_AND_wci_wReset_n_8_336__ETC___d3423 ;

  // rule RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_T
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_T =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd8 &&
	     cpReq[61:60] == 2'd1 &&
	     cpReq[19:9] == 11'd0 &&
	     !wci_busy_8 &&
	     wci_respF_8$FULL_N &&
	     !dispatched ;

  // rule RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_F_F_T
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_F_F_T =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd8 &&
	     cpReq[61:60] != 2'd2 &&
	     (cpReq[61:60] != 2'd1 || cpReq[19:9] != 11'd0) &&
	     cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_AND_NOT_w_ETC___d3460 ;

  // rule RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_F_F_F
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_F_F_F =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd8 &&
	     cpReq[61:60] != 2'd2 &&
	     (cpReq[61:60] != 2'd1 || cpReq[19:9] != 11'd0) &&
	     cpReq[9:6] != 4'h9 &&
	     NOT_cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_961_A_ETC___d3466 ;

  // rule RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_T_F
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_T_F =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd9 &&
	     cpReq[61:60] == 2'd2 &&
	     !wci_wReset_n_9 &&
	     NOT_wci_busy_9_496_473_AND_wci_wReset_n_9_476__ETC___d3486 ;

  // rule RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_T
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_T =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd9 &&
	     cpReq[61:60] == 2'd1 &&
	     cpReq[19:9] == 11'd0 &&
	     !wci_busy_9 &&
	     wci_respF_9$FULL_N &&
	     !dispatched ;

  // rule RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_F_F_T
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_F_F_T =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd9 &&
	     cpReq[61:60] != 2'd2 &&
	     (cpReq[61:60] != 2'd1 || cpReq[19:9] != 11'd0) &&
	     cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_AND_NOT_w_ETC___d3523 ;

  // rule RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_F_F_F
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_F_F_F =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd9 &&
	     cpReq[61:60] != 2'd2 &&
	     (cpReq[61:60] != 2'd1 || cpReq[19:9] != 11'd0) &&
	     cpReq[9:6] != 4'h9 &&
	     NOT_cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_961_A_ETC___d3529 ;

  // rule RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_T_F
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_T_F =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd10 &&
	     cpReq[61:60] == 2'd2 &&
	     !wci_wReset_n_10 &&
	     NOT_wci_busy_10_636_536_AND_wci_wReset_n_10_61_ETC___d3549 ;

  // rule RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_T
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_T =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd10 &&
	     cpReq[61:60] == 2'd1 &&
	     cpReq[19:9] == 11'd0 &&
	     !wci_busy_10 &&
	     wci_respF_10$FULL_N &&
	     !dispatched ;

  // rule RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd10 &&
	     cpReq[61:60] != 2'd2 &&
	     (cpReq[61:60] != 2'd1 || cpReq[19:9] != 11'd0) &&
	     cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_AND_NOT_w_ETC___d3586 ;

  // rule RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd10 &&
	     cpReq[61:60] != 2'd2 &&
	     (cpReq[61:60] != 2'd1 || cpReq[19:9] != 11'd0) &&
	     cpReq[9:6] != 4'h9 &&
	     NOT_cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_961_A_ETC___d3592 ;

  // rule RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_T_F
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_T_F =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd11 &&
	     cpReq[61:60] == 2'd2 &&
	     !wci_wReset_n_11 &&
	     NOT_wci_busy_11_776_599_AND_wci_wReset_n_11_75_ETC___d3612 ;

  // rule RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_T
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_T =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd11 &&
	     cpReq[61:60] == 2'd1 &&
	     cpReq[19:9] == 11'd0 &&
	     !wci_busy_11 &&
	     wci_respF_11$FULL_N &&
	     !dispatched ;

  // rule RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd11 &&
	     cpReq[61:60] != 2'd2 &&
	     (cpReq[61:60] != 2'd1 || cpReq[19:9] != 11'd0) &&
	     cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_AND_NOT_w_ETC___d3649 ;

  // rule RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd11 &&
	     cpReq[61:60] != 2'd2 &&
	     (cpReq[61:60] != 2'd1 || cpReq[19:9] != 11'd0) &&
	     cpReq[9:6] != 4'h9 &&
	     NOT_cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_961_A_ETC___d3655 ;

  // rule RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd12 &&
	     cpReq[61:60] == 2'd2 &&
	     !wci_wReset_n_12 &&
	     NOT_wci_busy_12_916_662_AND_wci_wReset_n_12_89_ETC___d3675 ;

  // rule RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd12 &&
	     cpReq[61:60] == 2'd1 &&
	     cpReq[19:9] == 11'd0 &&
	     !wci_busy_12 &&
	     wci_respF_12$FULL_N &&
	     !dispatched ;

  // rule RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd12 &&
	     cpReq[61:60] != 2'd2 &&
	     (cpReq[61:60] != 2'd1 || cpReq[19:9] != 11'd0) &&
	     cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_AND_NOT_w_ETC___d3712 ;

  // rule RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd12 &&
	     cpReq[61:60] != 2'd2 &&
	     (cpReq[61:60] != 2'd1 || cpReq[19:9] != 11'd0) &&
	     cpReq[9:6] != 4'h9 &&
	     NOT_cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_961_A_ETC___d3718 ;

  // rule RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd13 &&
	     cpReq[61:60] == 2'd2 &&
	     !wci_wReset_n_13 &&
	     NOT_wci_busy_13_056_725_AND_wci_wReset_n_13_03_ETC___d3738 ;

  // rule RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd13 &&
	     cpReq[61:60] == 2'd1 &&
	     cpReq[19:9] == 11'd0 &&
	     !wci_busy_13 &&
	     wci_respF_13$FULL_N &&
	     !dispatched ;

  // rule RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd13 &&
	     cpReq[61:60] != 2'd2 &&
	     (cpReq[61:60] != 2'd1 || cpReq[19:9] != 11'd0) &&
	     cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_AND_NOT_w_ETC___d3775 ;

  // rule RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd13 &&
	     cpReq[61:60] != 2'd2 &&
	     (cpReq[61:60] != 2'd1 || cpReq[19:9] != 11'd0) &&
	     cpReq[9:6] != 4'h9 &&
	     NOT_cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_961_A_ETC___d3781 ;

  // rule RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd14 &&
	     cpReq[61:60] == 2'd2 &&
	     !wci_wReset_n_14 &&
	     NOT_wci_busy_14_196_788_AND_wci_wReset_n_14_17_ETC___d3801 ;

  // rule RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd14 &&
	     cpReq[61:60] == 2'd1 &&
	     cpReq[19:9] == 11'd0 &&
	     !wci_busy_14 &&
	     wci_respF_14$FULL_N &&
	     !dispatched ;

  // rule RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd14 &&
	     cpReq[61:60] != 2'd2 &&
	     (cpReq[61:60] != 2'd1 || cpReq[19:9] != 11'd0) &&
	     cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_AND_NOT_w_ETC___d3838 ;

  // rule RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd14 &&
	     cpReq[61:60] != 2'd2 &&
	     (cpReq[61:60] != 2'd1 || cpReq[19:9] != 11'd0) &&
	     cpReq[9:6] != 4'h9 &&
	     NOT_cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_961_A_ETC___d3844 ;

  // rule RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 != 4'd0 &&
	     _theResult_____1__h76796 != 4'd1 &&
	     _theResult_____1__h76796 != 4'd2 &&
	     _theResult_____1__h76796 != 4'd3 &&
	     _theResult_____1__h76796 != 4'd4 &&
	     _theResult_____1__h76796 != 4'd5 &&
	     _theResult_____1__h76796 != 4'd6 &&
	     _theResult_____1__h76796 != 4'd7 &&
	     _theResult_____1__h76796 != 4'd8 &&
	     _theResult_____1__h76796 != 4'd9 &&
	     _theResult_____1__h76796 != 4'd10 &&
	     _theResult_____1__h76796 != 4'd11 &&
	     _theResult_____1__h76796 != 4'd12 &&
	     _theResult_____1__h76796 != 4'd13 &&
	     _theResult_____1__h76796 != 4'd14 &&
	     !dispatched ;

  // rule RL_cpDispatch_F_F_F_T
  assign WILL_FIRE_RL_cpDispatch_F_F_F_T =
	     cpReq[64:62] == 3'd0 && !dispatched ;

  // rule RL_cpDispatch_F_F_F_F_T_T_F
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_T_T_F =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     _theResult_____1__h76814 == 4'd0 &&
	     cpReq[37:36] == 2'd2 &&
	     !wci_wReset_n &&
	     NOT_wci_busy_36_886_AND_wci_wReset_n_16_OR_wci_ETC___d2904 ;

  // rule RL_cpDispatch_F_F_F_F_T_F_T_F
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_T_F_T_F =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     _theResult_____1__h76814 == 4'd0 &&
	     cpReq[37:36] == 2'd1 &&
	     cpReq[19:9] == 11'd0 &&
	     !wci_wReset_n &&
	     NOT_wci_busy_36_886_AND_wci_wReset_n_16_OR_wci_ETC___d2904 ;

  // rule RL_cpDispatch_F_F_F_F_T_F_F_T
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_T_F_F_T =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d3932 ;

  // rule RL_cpDispatch_F_F_F_F_T_F_F_F_T
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_T_F_F_F_T =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d3941 ;

  // rule RL_cpDispatch_F_F_F_F_T_F_F_F_F_T
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_T_F_F_F_F_T =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d3951 ;

  // rule RL_cpDispatch_F_F_F_F_T_F_F_F_F_F_T
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_T_F_F_F_F_F_T =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     _theResult_____1__h76814 == 4'd0 &&
	     cpReq[37:36] != 2'd2 &&
	     (cpReq[37:36] != 2'd1 || cpReq[19:9] != 11'd0) &&
	     cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_AND_NOT_w_ETC___d2953 ;

  // rule RL_cpDispatch_F_F_F_F_T_F_F_F_F_F_F
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_T_F_F_F_F_F_F =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     NOT_cpReq_363_BITS_64_TO_62_364_EQ_3_877_885_A_ETC___d3976 ;

  // rule RL_cpDispatch_F_F_F_F_F_T_T_F
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_T_F =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     _theResult_____1__h76814 == 4'd1 &&
	     cpReq[37:36] == 2'd2 &&
	     !wci_wReset_n_1 &&
	     NOT_wci_busy_1_76_969_AND_wci_wReset_n_1_56_OR_ETC___d2982 ;

  // rule RL_cpDispatch_F_F_F_F_F_T_F_T_F
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_F_T_F =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     _theResult_____1__h76814 == 4'd1 &&
	     cpReq[37:36] == 2'd1 &&
	     cpReq[19:9] == 11'd0 &&
	     !wci_wReset_n_1 &&
	     NOT_wci_busy_1_76_969_AND_wci_wReset_n_1_56_OR_ETC___d2982 ;

  // rule RL_cpDispatch_F_F_F_F_F_T_F_F_T
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_F_F_T =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4010 ;

  // rule RL_cpDispatch_F_F_F_F_F_T_F_F_F_T
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_F_F_F_T =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4019 ;

  // rule RL_cpDispatch_F_F_F_F_F_T_F_F_F_F_T
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_F_F_F_F_T =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4029 ;

  // rule RL_cpDispatch_F_F_F_F_F_T_F_F_F_F_F_T
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_F_F_F_F_F_T =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     _theResult_____1__h76814 == 4'd1 &&
	     cpReq[37:36] != 2'd2 &&
	     (cpReq[37:36] != 2'd1 || cpReq[19:9] != 11'd0) &&
	     cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_AND_NOT_w_ETC___d3019 ;

  // rule RL_cpDispatch_F_F_F_F_F_T_F_F_F_F_F_F
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_F_F_F_F_F_F =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     NOT_cpReq_363_BITS_64_TO_62_364_EQ_3_877_885_A_ETC___d4052 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_T_T_F
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_T_F =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     _theResult_____1__h76814 == 4'd2 &&
	     cpReq[37:36] == 2'd2 &&
	     !wci_wReset_n_2 &&
	     NOT_wci_busy_2_16_032_AND_wci_wReset_n_2_96_OR_ETC___d3045 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_T_F_T_F
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_F_T_F =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     _theResult_____1__h76814 == 4'd2 &&
	     cpReq[37:36] == 2'd1 &&
	     cpReq[19:9] == 11'd0 &&
	     !wci_wReset_n_2 &&
	     NOT_wci_busy_2_16_032_AND_wci_wReset_n_2_96_OR_ETC___d3045 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_T_F_F_T
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_F_F_T =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4086 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_T_F_F_F_T
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_F_F_F_T =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4095 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_T_F_F_F_F_T
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_F_F_F_F_T =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4105 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_T_F_F_F_F_F_T
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_F_F_F_F_F_T =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     _theResult_____1__h76814 == 4'd2 &&
	     cpReq[37:36] != 2'd2 &&
	     (cpReq[37:36] != 2'd1 || cpReq[19:9] != 11'd0) &&
	     cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_AND_NOT_w_ETC___d3082 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_T_F_F_F_F_F_F
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_F_F_F_F_F_F =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     NOT_cpReq_363_BITS_64_TO_62_364_EQ_3_877_885_A_ETC___d4128 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_T_T_F
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_T_F =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     _theResult_____1__h76814 == 4'd3 &&
	     cpReq[37:36] == 2'd2 &&
	     !wci_wReset_n_3 &&
	     NOT_wci_busy_3_56_095_AND_wci_wReset_n_3_36_OR_ETC___d3108 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_T_F_T_F
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_F_T_F =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     _theResult_____1__h76814 == 4'd3 &&
	     cpReq[37:36] == 2'd1 &&
	     cpReq[19:9] == 11'd0 &&
	     !wci_wReset_n_3 &&
	     NOT_wci_busy_3_56_095_AND_wci_wReset_n_3_36_OR_ETC___d3108 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_T_F_F_T
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_F_F_T =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4162 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_T_F_F_F_T
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_F_F_F_T =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4171 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_T_F_F_F_F_T
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_F_F_F_F_T =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4181 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_T_F_F_F_F_F_T
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_F_F_F_F_F_T =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     _theResult_____1__h76814 == 4'd3 &&
	     cpReq[37:36] != 2'd2 &&
	     (cpReq[37:36] != 2'd1 || cpReq[19:9] != 11'd0) &&
	     cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_AND_NOT_w_ETC___d3145 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_T_F_F_F_F_F_F
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_F_F_F_F_F_F =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     NOT_cpReq_363_BITS_64_TO_62_364_EQ_3_877_885_A_ETC___d4204 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_F_T_T_F
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_T_F =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     _theResult_____1__h76814 == 4'd4 &&
	     cpReq[37:36] == 2'd2 &&
	     !wci_wReset_n_4 &&
	     NOT_wci_busy_4_96_158_AND_wci_wReset_n_4_76_OR_ETC___d3171 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_F_T_F_T_F
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_F_T_F =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     _theResult_____1__h76814 == 4'd4 &&
	     cpReq[37:36] == 2'd1 &&
	     cpReq[19:9] == 11'd0 &&
	     !wci_wReset_n_4 &&
	     NOT_wci_busy_4_96_158_AND_wci_wReset_n_4_76_OR_ETC___d3171 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_F_T_F_F_T
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_F_F_T =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4238 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_F_T_F_F_F_T
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_F_F_F_T =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4247 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_F_T_F_F_F_F_T
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_F_F_F_F_T =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4257 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     _theResult_____1__h76814 == 4'd4 &&
	     cpReq[37:36] != 2'd2 &&
	     (cpReq[37:36] != 2'd1 || cpReq[19:9] != 11'd0) &&
	     cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_AND_NOT_w_ETC___d3208 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     NOT_cpReq_363_BITS_64_TO_62_364_EQ_3_877_885_A_ETC___d4280 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_T_F
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_T_F =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     _theResult_____1__h76814 == 4'd5 &&
	     cpReq[37:36] == 2'd2 &&
	     !wci_wReset_n_5 &&
	     NOT_wci_busy_5_36_221_AND_wci_wReset_n_5_16_OR_ETC___d3234 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_F_T_F
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_F_T_F =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     _theResult_____1__h76814 == 4'd5 &&
	     cpReq[37:36] == 2'd1 &&
	     cpReq[19:9] == 11'd0 &&
	     !wci_wReset_n_5 &&
	     NOT_wci_busy_5_36_221_AND_wci_wReset_n_5_16_OR_ETC___d3234 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_F_F_T
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_F_F_T =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4314 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_F_F_F_T
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_F_F_F_T =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4323 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4333 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     _theResult_____1__h76814 == 4'd5 &&
	     cpReq[37:36] != 2'd2 &&
	     (cpReq[37:36] != 2'd1 || cpReq[19:9] != 11'd0) &&
	     cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_AND_NOT_w_ETC___d3271 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     NOT_cpReq_363_BITS_64_TO_62_364_EQ_3_877_885_A_ETC___d4356 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_T_F
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_T_F =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     _theResult_____1__h76814 == 4'd6 &&
	     cpReq[37:36] == 2'd2 &&
	     !wci_wReset_n_6 &&
	     NOT_wci_busy_6_076_284_AND_wci_wReset_n_6_056__ETC___d3297 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_F_T_F
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_F_T_F =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     _theResult_____1__h76814 == 4'd6 &&
	     cpReq[37:36] == 2'd1 &&
	     cpReq[19:9] == 11'd0 &&
	     !wci_wReset_n_6 &&
	     NOT_wci_busy_6_076_284_AND_wci_wReset_n_6_056__ETC___d3297 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_F_F_T
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_F_F_T =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4390 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4399 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4409 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     _theResult_____1__h76814 == 4'd6 &&
	     cpReq[37:36] != 2'd2 &&
	     (cpReq[37:36] != 2'd1 || cpReq[19:9] != 11'd0) &&
	     cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_AND_NOT_w_ETC___d3334 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     NOT_cpReq_363_BITS_64_TO_62_364_EQ_3_877_885_A_ETC___d4432 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_T_F
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_T_F =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     _theResult_____1__h76814 == 4'd7 &&
	     cpReq[37:36] == 2'd2 &&
	     !wci_wReset_n_7 &&
	     NOT_wci_busy_7_216_347_AND_wci_wReset_n_7_196__ETC___d3360 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     _theResult_____1__h76814 == 4'd7 &&
	     cpReq[37:36] == 2'd1 &&
	     cpReq[19:9] == 11'd0 &&
	     !wci_wReset_n_7 &&
	     NOT_wci_busy_7_216_347_AND_wci_wReset_n_7_196__ETC___d3360 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4466 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4475 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4485 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     _theResult_____1__h76814 == 4'd7 &&
	     cpReq[37:36] != 2'd2 &&
	     (cpReq[37:36] != 2'd1 || cpReq[19:9] != 11'd0) &&
	     cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_AND_NOT_w_ETC___d3397 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     NOT_cpReq_363_BITS_64_TO_62_364_EQ_3_877_885_A_ETC___d4508 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     _theResult_____1__h76814 == 4'd8 &&
	     cpReq[37:36] == 2'd2 &&
	     !wci_wReset_n_8 &&
	     NOT_wci_busy_8_356_410_AND_wci_wReset_n_8_336__ETC___d3423 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     _theResult_____1__h76814 == 4'd8 &&
	     cpReq[37:36] == 2'd1 &&
	     cpReq[19:9] == 11'd0 &&
	     !wci_wReset_n_8 &&
	     NOT_wci_busy_8_356_410_AND_wci_wReset_n_8_336__ETC___d3423 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4542 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4551 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4561 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     _theResult_____1__h76814 == 4'd8 &&
	     cpReq[37:36] != 2'd2 &&
	     (cpReq[37:36] != 2'd1 || cpReq[19:9] != 11'd0) &&
	     cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_AND_NOT_w_ETC___d3460 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     NOT_cpReq_363_BITS_64_TO_62_364_EQ_3_877_885_A_ETC___d4584 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     _theResult_____1__h76814 == 4'd9 &&
	     cpReq[37:36] == 2'd2 &&
	     !wci_wReset_n_9 &&
	     NOT_wci_busy_9_496_473_AND_wci_wReset_n_9_476__ETC___d3486 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     _theResult_____1__h76814 == 4'd9 &&
	     cpReq[37:36] == 2'd1 &&
	     cpReq[19:9] == 11'd0 &&
	     !wci_wReset_n_9 &&
	     NOT_wci_busy_9_496_473_AND_wci_wReset_n_9_476__ETC___d3486 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4618 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4627 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4637 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     _theResult_____1__h76814 == 4'd9 &&
	     cpReq[37:36] != 2'd2 &&
	     (cpReq[37:36] != 2'd1 || cpReq[19:9] != 11'd0) &&
	     cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_AND_NOT_w_ETC___d3523 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     NOT_cpReq_363_BITS_64_TO_62_364_EQ_3_877_885_A_ETC___d4660 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     _theResult_____1__h76814 == 4'd10 &&
	     cpReq[37:36] == 2'd2 &&
	     !wci_wReset_n_10 &&
	     NOT_wci_busy_10_636_536_AND_wci_wReset_n_10_61_ETC___d3549 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     _theResult_____1__h76814 == 4'd10 &&
	     cpReq[37:36] == 2'd1 &&
	     cpReq[19:9] == 11'd0 &&
	     !wci_wReset_n_10 &&
	     NOT_wci_busy_10_636_536_AND_wci_wReset_n_10_61_ETC___d3549 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4694 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4703 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4713 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     _theResult_____1__h76814 == 4'd10 &&
	     cpReq[37:36] != 2'd2 &&
	     (cpReq[37:36] != 2'd1 || cpReq[19:9] != 11'd0) &&
	     cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_AND_NOT_w_ETC___d3586 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     NOT_cpReq_363_BITS_64_TO_62_364_EQ_3_877_885_A_ETC___d4736 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     _theResult_____1__h76814 == 4'd11 &&
	     cpReq[37:36] == 2'd2 &&
	     !wci_wReset_n_11 &&
	     NOT_wci_busy_11_776_599_AND_wci_wReset_n_11_75_ETC___d3612 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     _theResult_____1__h76814 == 4'd11 &&
	     cpReq[37:36] == 2'd1 &&
	     cpReq[19:9] == 11'd0 &&
	     !wci_wReset_n_11 &&
	     NOT_wci_busy_11_776_599_AND_wci_wReset_n_11_75_ETC___d3612 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4770 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4779 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4789 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     _theResult_____1__h76814 == 4'd11 &&
	     cpReq[37:36] != 2'd2 &&
	     (cpReq[37:36] != 2'd1 || cpReq[19:9] != 11'd0) &&
	     cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_AND_NOT_w_ETC___d3649 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     NOT_cpReq_363_BITS_64_TO_62_364_EQ_3_877_885_A_ETC___d4812 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     _theResult_____1__h76814 == 4'd12 &&
	     cpReq[37:36] == 2'd2 &&
	     !wci_wReset_n_12 &&
	     NOT_wci_busy_12_916_662_AND_wci_wReset_n_12_89_ETC___d3675 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     _theResult_____1__h76814 == 4'd12 &&
	     cpReq[37:36] == 2'd1 &&
	     cpReq[19:9] == 11'd0 &&
	     !wci_wReset_n_12 &&
	     NOT_wci_busy_12_916_662_AND_wci_wReset_n_12_89_ETC___d3675 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4846 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4855 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4865 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     _theResult_____1__h76814 == 4'd12 &&
	     cpReq[37:36] != 2'd2 &&
	     (cpReq[37:36] != 2'd1 || cpReq[19:9] != 11'd0) &&
	     cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_AND_NOT_w_ETC___d3712 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     NOT_cpReq_363_BITS_64_TO_62_364_EQ_3_877_885_A_ETC___d4888 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     _theResult_____1__h76814 == 4'd13 &&
	     cpReq[37:36] == 2'd2 &&
	     !wci_wReset_n_13 &&
	     NOT_wci_busy_13_056_725_AND_wci_wReset_n_13_03_ETC___d3738 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     _theResult_____1__h76814 == 4'd13 &&
	     cpReq[37:36] == 2'd1 &&
	     cpReq[19:9] == 11'd0 &&
	     !wci_wReset_n_13 &&
	     NOT_wci_busy_13_056_725_AND_wci_wReset_n_13_03_ETC___d3738 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4922 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4931 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4941 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     _theResult_____1__h76814 == 4'd13 &&
	     cpReq[37:36] != 2'd2 &&
	     (cpReq[37:36] != 2'd1 || cpReq[19:9] != 11'd0) &&
	     cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_AND_NOT_w_ETC___d3775 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     NOT_cpReq_363_BITS_64_TO_62_364_EQ_3_877_885_A_ETC___d4964 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     _theResult_____1__h76814 == 4'd14 &&
	     cpReq[37:36] == 2'd2 &&
	     !wci_wReset_n_14 &&
	     NOT_wci_busy_14_196_788_AND_wci_wReset_n_14_17_ETC___d3801 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     _theResult_____1__h76814 == 4'd14 &&
	     cpReq[37:36] == 2'd1 &&
	     cpReq[19:9] == 11'd0 &&
	     !wci_wReset_n_14 &&
	     NOT_wci_busy_14_196_788_AND_wci_wReset_n_14_17_ETC___d3801 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4998 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d5007 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d5017 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     _theResult_____1__h76814 == 4'd14 &&
	     cpReq[37:36] != 2'd2 &&
	     (cpReq[37:36] != 2'd1 || cpReq[19:9] != 11'd0) &&
	     cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_AND_NOT_w_ETC___d3838 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     NOT_cpReq_363_BITS_64_TO_62_364_EQ_3_877_885_A_ETC___d5040 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     NOT_cpReq_363_BITS_64_TO_62_364_EQ_0_881_886_A_ETC___d5073 ;

  // rule RL_completeWorkerWrite
  assign WILL_FIRE_RL_completeWorkerWrite =
	     IF_wrkAct_077_EQ_0_078_THEN_wci_respF_i_notEmp_ETC___d6132 &&
	     cpReq[64:62] == 3'd3 &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_F &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_F &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_F &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_F &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_F &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_F &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_F &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_F &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_T_F &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_T_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_F &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_F &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_T_F &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_T_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_F_F_F &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_F_F_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_F_T_F_F &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_F_T_F_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_F_T_T_F &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_T_F &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_T_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_F_F_F &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_F_F_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_F_T_F_F &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_F_T_F_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_F_T_T_F &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_F_T_T_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_T_F &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_T_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_F_F_F &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_F_F_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_F_T_F_F &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_F_T_F_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_F_T_T_F &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_F_T_T_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_T_F &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_T_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_F_F_F &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_F_F_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_F_T_F_F &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_F_T_F_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_F_T_T_F &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_F_T_T_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_T_F &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_T_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_F_F_F &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_F_T_F_F &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_F_F_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_F_T_F_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_F_T_T_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_F_T_T_F &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_T_F &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_T_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_F_F_F_F &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_F_F_F_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_F_F_T_F_F &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_F_F_T_F_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_F_F_T_T_F &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_F_F_T_T_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_T_F &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_F_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_T_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_F_F_F_F &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_F_F_F_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_F_F_T_F_F &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_F_F_T_F_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_F_F_T_T_F &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_F_F_T_T_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_F_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_T_F &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_T_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_F_F_F_F &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_F_F_F_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_F_F_T_F_F &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_F_F_T_F_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_F_F_T_T_F &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_F_F_T_T_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_F_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_T_F &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_T_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_T_F_F_F_F &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_T_F_F_F_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_T_F_F_T_F_F &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_T_F_F_T_F_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_T_F_F_T_T_F &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_T_F_F_T_T_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_T_F_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_T_T_F &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_F_T_T_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_T_F_F_F_F &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_T_F_F_T_F_F &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_T_F_F_T_F_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_T_F_F_T_T_F &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_T_F_F_F_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_T_F_F_T_T_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_T_F_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_T_T_F &&
	     !WILL_FIRE_RL_cpDispatch_F_F_T_T_T_T ;

  // rule RL_completeWorkerRead
  assign WILL_FIRE_RL_completeWorkerRead =
	     cpRespF$FULL_N &&
	     IF_wrkAct_077_EQ_0_078_THEN_wci_respF_i_notEmp_ETC___d6132 &&
	     cpReq[64:62] != 3'd0 &&
	     cpReq[64:62] != 3'd1 &&
	     cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_T_F &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_T_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_F_F_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_F_T_F &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_F_T_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_T_F &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_T_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_F_F_F_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_F_F_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_F_T_F &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_F_T_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_T_F &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_T_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_F_F_F_F_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_F_F_F_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_F_F_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_F_T_F &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_F_T_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_T_F &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_T_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_F_F_F_F_F_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_F_F_F_F_F_F &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_F_F_F_F_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_F_F_F_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_F_F_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_F_T_F &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_F_T_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_T_F &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_T_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_F_F_F_F_F_F &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_F_F_F_F_F_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_F_F_F_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_F_F_F_F_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_F_F_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_F_T_F &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_F_T_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_T_F &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_T_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_F_F_F_F_F_F &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_F_F_F_F_F_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_F_F_F_F_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_F_F_F_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_F_F_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_F_T_F &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_F_T_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_T_F &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_T_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_T_F_F_F_F_F_F &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_T_F_F_F_F_F_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_T_F_F_F_F_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_T_F_F_F_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_T_F_F_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_T_F_T_T &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_T_F_T_F &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_T_T_F &&
	     !WILL_FIRE_RL_cpDispatch_F_F_F_F_T_T_T &&
	     !WILL_FIRE_RL_responseAdminRd ;

  // rule RL_reqRcv
  assign WILL_FIRE_RL_reqRcv = cpReqF$EMPTY_N && cpReq[64:62] == 3'd0 ;

  // rule RL_cpDispatch_T_F_F_F_F_T_T
  assign WILL_FIRE_RL_cpDispatch_T_F_F_F_F_T_T =
	     cpReq[64:62] == 3'd1 && cpReq[11:4] == 8'h34 && cpReq[59] &&
	     !dispatched ;

  // rule RL_cpDispatch_T_F_F_F_F_T_F
  assign WILL_FIRE_RL_cpDispatch_T_F_F_F_F_T_F =
	     cpReq[64:62] == 3'd1 && cpReq[11:4] == 8'h34 && !cpReq[59] &&
	     !dispatched ;

`ifdef not
  // rule RL_rom_serverAdapter_stageReadResponseAlways
  assign WILL_FIRE_RL_rom_serverAdapter_stageReadResponseAlways =
	     CAN_FIRE_RL_cpDispatch_F_T_F_F && !WILL_FIRE_RL_responseAdminRd ;

  // rule RL_rom_serverAdapter_outData_enqAndDeq
  assign WILL_FIRE_RL_rom_serverAdapter_outData_enqAndDeq =
	     rom_serverAdapter_outDataCore$EMPTY_N &&
	     rom_serverAdapter_outDataCore$FULL_N &&
	     rom_serverAdapter_outData_deqCalled$whas &&
	     rom_serverAdapter_outData_enqData$whas ;
`endif
	      
  // rule RL_cpDispatch_F_F_T_T_F_F_T_T_F
  assign WILL_FIRE_RL_cpDispatch_F_F_T_T_F_F_T_T_F =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd0 &&
	     cpReq[61:60] != 2'd2 &&
	     cpReq[9:6] == 4'h9 &&
	     cpReq[37] &&
	     NOT_cpReq_363_BIT_36_924_932_AND_NOT_wci_busy__ETC___d2933 ;

  // rule RL_cpDispatch_F_F_T_T_F_F_T_F_F
  assign WILL_FIRE_RL_cpDispatch_F_F_T_T_F_F_T_F_F =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd0 &&
	     cpReq[61:60] != 2'd2 &&
	     cpReq[9:6] == 4'h9 &&
	     !cpReq[37] &&
	     NOT_cpReq_363_BIT_36_924_932_AND_NOT_wci_busy__ETC___d2933 ;

  // rule RL_cpDispatch_F_F_T_T_T_T
  assign WILL_FIRE_RL_cpDispatch_F_F_T_T_T_T =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd0 &&
	     cpReq[61:60] == 2'd2 &&
	     wci_wReset_n_16_AND_NOT_wci_busy_36_886_AND_NO_ETC___d2889 ;

  // rule RL_cpDispatch_F_F_T_T_F_F_T_T_T
  assign WILL_FIRE_RL_cpDispatch_F_F_T_T_F_F_T_T_T =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd0 &&
	     cpReq[61:60] != 2'd2 &&
	     cpReq[9:6] == 4'h9 &&
	     cpReq[37] &&
	     cpReq_363_BIT_36_924_AND_NOT_wci_busy_36_886_A_ETC___d2925 ;

  // rule RL_cpDispatch_F_F_T_T_F_F_T_F_T
  assign WILL_FIRE_RL_cpDispatch_F_F_T_T_F_F_T_F_T =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd0 &&
	     cpReq[61:60] != 2'd2 &&
	     cpReq[9:6] == 4'h9 &&
	     !cpReq[37] &&
	     cpReq_363_BIT_36_924_AND_NOT_wci_busy_36_886_A_ETC___d2925 ;

  // rule RL_cpDispatch_F_F_F_F_T_T_T
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_T_T_T =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     _theResult_____1__h76814 == 4'd0 &&
	     cpReq[37:36] == 2'd2 &&
	     wci_wReset_n_16_AND_NOT_wci_busy_36_886_AND_NO_ETC___d2889 ;

  // rule RL_cpDispatch_F_F_F_F_T_F_T_T
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_T_F_T_T =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     _theResult_____1__h76814 == 4'd0 &&
	     cpReq[37:36] == 2'd1 &&
	     cpReq[19:9] == 11'd0 &&
	     wci_wReset_n_16_AND_NOT_wci_busy_36_886_AND_NO_ETC___d2889 ;

  // rule RL_cpDispatch_F_F_T_F_T_F_F_T_T_F
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_T_F_F_T_T_F =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd1 &&
	     cpReq[61:60] != 2'd2 &&
	     cpReq[9:6] == 4'h9 &&
	     cpReq[37] &&
	     NOT_cpReq_363_BIT_36_924_932_AND_NOT_wci_busy__ETC___d3000 ;

  // rule RL_cpDispatch_F_F_T_F_T_F_F_T_F_F
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_T_F_F_T_F_F =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd1 &&
	     cpReq[61:60] != 2'd2 &&
	     cpReq[9:6] == 4'h9 &&
	     !cpReq[37] &&
	     NOT_cpReq_363_BIT_36_924_932_AND_NOT_wci_busy__ETC___d3000 ;

  // rule RL_cpDispatch_F_F_T_F_T_T_T
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_T_T_T =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd1 &&
	     cpReq[61:60] == 2'd2 &&
	     wci_wReset_n_1_56_AND_NOT_wci_busy_1_76_969_AN_ETC___d2972 ;

  // rule RL_cpDispatch_F_F_T_F_T_F_F_T_T_T
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_T_F_F_T_T_T =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd1 &&
	     cpReq[61:60] != 2'd2 &&
	     cpReq[9:6] == 4'h9 &&
	     cpReq[37] &&
	     cpReq_363_BIT_36_924_AND_NOT_wci_busy_1_76_969_ETC___d2993 ;

  // rule RL_cpDispatch_F_F_T_F_T_F_F_T_F_T
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_T_F_F_T_F_T =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd1 &&
	     cpReq[61:60] != 2'd2 &&
	     cpReq[9:6] == 4'h9 &&
	     !cpReq[37] &&
	     cpReq_363_BIT_36_924_AND_NOT_wci_busy_1_76_969_ETC___d2993 ;

  // rule RL_cpDispatch_F_F_F_F_F_T_T_T
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_T_T =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     _theResult_____1__h76814 == 4'd1 &&
	     cpReq[37:36] == 2'd2 &&
	     wci_wReset_n_1_56_AND_NOT_wci_busy_1_76_969_AN_ETC___d2972 ;

  // rule RL_cpDispatch_F_F_F_F_F_T_F_T_T
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_F_T_T =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     _theResult_____1__h76814 == 4'd1 &&
	     cpReq[37:36] == 2'd1 &&
	     cpReq[19:9] == 11'd0 &&
	     wci_wReset_n_1_56_AND_NOT_wci_busy_1_76_969_AN_ETC___d2972 ;

  // rule RL_cpDispatch_F_F_T_F_F_T_F_F_T_T_F
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_F_F_T_T_F =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd2 &&
	     cpReq[61:60] != 2'd2 &&
	     cpReq[9:6] == 4'h9 &&
	     cpReq[37] &&
	     NOT_cpReq_363_BIT_36_924_932_AND_NOT_wci_busy__ETC___d3063 ;

  // rule RL_cpDispatch_F_F_T_F_F_T_F_F_T_F_F
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_F_F_T_F_F =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd2 &&
	     cpReq[61:60] != 2'd2 &&
	     cpReq[9:6] == 4'h9 &&
	     !cpReq[37] &&
	     NOT_cpReq_363_BIT_36_924_932_AND_NOT_wci_busy__ETC___d3063 ;

  // rule RL_cpDispatch_F_F_T_F_F_T_T_T
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_T_T =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd2 &&
	     cpReq[61:60] == 2'd2 &&
	     wci_wReset_n_2_96_AND_NOT_wci_busy_2_16_032_AN_ETC___d3035 ;

  // rule RL_cpDispatch_F_F_T_F_F_T_F_F_T_T_T
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_F_F_T_T_T =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd2 &&
	     cpReq[61:60] != 2'd2 &&
	     cpReq[9:6] == 4'h9 &&
	     cpReq[37] &&
	     cpReq_363_BIT_36_924_AND_NOT_wci_busy_2_16_032_ETC___d3056 ;

  // rule RL_cpDispatch_F_F_T_F_F_T_F_F_T_F_T
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_F_F_T_F_T =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd2 &&
	     cpReq[61:60] != 2'd2 &&
	     cpReq[9:6] == 4'h9 &&
	     !cpReq[37] &&
	     cpReq_363_BIT_36_924_AND_NOT_wci_busy_2_16_032_ETC___d3056 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_T_T_T
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_T_T =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     _theResult_____1__h76814 == 4'd2 &&
	     cpReq[37:36] == 2'd2 &&
	     wci_wReset_n_2_96_AND_NOT_wci_busy_2_16_032_AN_ETC___d3035 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_T_F_T_T
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_F_T_T =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     _theResult_____1__h76814 == 4'd2 &&
	     cpReq[37:36] == 2'd1 &&
	     cpReq[19:9] == 11'd0 &&
	     wci_wReset_n_2_96_AND_NOT_wci_busy_2_16_032_AN_ETC___d3035 ;

  // rule RL_cpDispatch_F_F_T_F_F_F_T_F_F_T_T_F
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_F_F_T_T_F =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd3 &&
	     cpReq[61:60] != 2'd2 &&
	     cpReq[9:6] == 4'h9 &&
	     cpReq[37] &&
	     NOT_cpReq_363_BIT_36_924_932_AND_NOT_wci_busy__ETC___d3126 ;

  // rule RL_cpDispatch_F_F_T_F_F_F_T_F_F_T_F_F
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_F_F_T_F_F =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd3 &&
	     cpReq[61:60] != 2'd2 &&
	     cpReq[9:6] == 4'h9 &&
	     !cpReq[37] &&
	     NOT_cpReq_363_BIT_36_924_932_AND_NOT_wci_busy__ETC___d3126 ;

  // rule RL_cpDispatch_F_F_T_F_F_F_T_T_T
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_T_T =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd3 &&
	     cpReq[61:60] == 2'd2 &&
	     wci_wReset_n_3_36_AND_NOT_wci_busy_3_56_095_AN_ETC___d3098 ;

  // rule RL_cpDispatch_F_F_T_F_F_F_T_F_F_T_T_T
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_F_F_T_T_T =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd3 &&
	     cpReq[61:60] != 2'd2 &&
	     cpReq[9:6] == 4'h9 &&
	     cpReq[37] &&
	     cpReq_363_BIT_36_924_AND_NOT_wci_busy_3_56_095_ETC___d3119 ;

  // rule RL_cpDispatch_F_F_T_F_F_F_T_F_F_T_F_T
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_F_F_T_F_T =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd3 &&
	     cpReq[61:60] != 2'd2 &&
	     cpReq[9:6] == 4'h9 &&
	     !cpReq[37] &&
	     cpReq_363_BIT_36_924_AND_NOT_wci_busy_3_56_095_ETC___d3119 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_T_T_T
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_T_T =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     _theResult_____1__h76814 == 4'd3 &&
	     cpReq[37:36] == 2'd2 &&
	     wci_wReset_n_3_36_AND_NOT_wci_busy_3_56_095_AN_ETC___d3098 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_T_F_T_T
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_F_T_T =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     _theResult_____1__h76814 == 4'd3 &&
	     cpReq[37:36] == 2'd1 &&
	     cpReq[19:9] == 11'd0 &&
	     wci_wReset_n_3_36_AND_NOT_wci_busy_3_56_095_AN_ETC___d3098 ;

  // rule RL_cpDispatch_F_F_T_F_F_F_F_T_F_F_T_T_F
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_F_F_T_T_F =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd4 &&
	     cpReq[61:60] != 2'd2 &&
	     cpReq[9:6] == 4'h9 &&
	     cpReq[37] &&
	     NOT_cpReq_363_BIT_36_924_932_AND_NOT_wci_busy__ETC___d3189 ;

  // rule RL_cpDispatch_F_F_T_F_F_F_F_T_F_F_T_F_F
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_F_F_T_F_F =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd4 &&
	     cpReq[61:60] != 2'd2 &&
	     cpReq[9:6] == 4'h9 &&
	     !cpReq[37] &&
	     NOT_cpReq_363_BIT_36_924_932_AND_NOT_wci_busy__ETC___d3189 ;

  // rule RL_cpDispatch_F_F_T_F_F_F_F_T_T_T
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_T_T =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd4 &&
	     cpReq[61:60] == 2'd2 &&
	     wci_wReset_n_4_76_AND_NOT_wci_busy_4_96_158_AN_ETC___d3161 ;

  // rule RL_cpDispatch_F_F_T_F_F_F_F_T_F_F_T_T_T
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_F_F_T_T_T =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd4 &&
	     cpReq[61:60] != 2'd2 &&
	     cpReq[9:6] == 4'h9 &&
	     cpReq[37] &&
	     cpReq_363_BIT_36_924_AND_NOT_wci_busy_4_96_158_ETC___d3182 ;

  // rule RL_cpDispatch_F_F_T_F_F_F_F_T_F_F_T_F_T
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_F_F_T_F_T =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd4 &&
	     cpReq[61:60] != 2'd2 &&
	     cpReq[9:6] == 4'h9 &&
	     !cpReq[37] &&
	     cpReq_363_BIT_36_924_AND_NOT_wci_busy_4_96_158_ETC___d3182 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_F_T_T_T
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_T_T =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     _theResult_____1__h76814 == 4'd4 &&
	     cpReq[37:36] == 2'd2 &&
	     wci_wReset_n_4_76_AND_NOT_wci_busy_4_96_158_AN_ETC___d3161 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_F_T_F_T_T
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_F_T_T =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     _theResult_____1__h76814 == 4'd4 &&
	     cpReq[37:36] == 2'd1 &&
	     cpReq[19:9] == 11'd0 &&
	     wci_wReset_n_4_76_AND_NOT_wci_busy_4_96_158_AN_ETC___d3161 ;

  // rule RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_F_T_T_F
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_F_T_T_F =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd5 &&
	     cpReq[61:60] != 2'd2 &&
	     cpReq[9:6] == 4'h9 &&
	     cpReq[37] &&
	     NOT_cpReq_363_BIT_36_924_932_AND_NOT_wci_busy__ETC___d3252 ;

  // rule RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_F_T_F_F
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_F_T_F_F =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd5 &&
	     cpReq[61:60] != 2'd2 &&
	     cpReq[9:6] == 4'h9 &&
	     !cpReq[37] &&
	     NOT_cpReq_363_BIT_36_924_932_AND_NOT_wci_busy__ETC___d3252 ;

  // rule RL_cpDispatch_F_F_T_F_F_F_F_F_T_T_T
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_T_T =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd5 &&
	     cpReq[61:60] == 2'd2 &&
	     wci_wReset_n_5_16_AND_NOT_wci_busy_5_36_221_AN_ETC___d3224 ;

  // rule RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_F_T_T_T
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_F_T_T_T =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd5 &&
	     cpReq[61:60] != 2'd2 &&
	     cpReq[9:6] == 4'h9 &&
	     cpReq[37] &&
	     cpReq_363_BIT_36_924_AND_NOT_wci_busy_5_36_221_ETC___d3245 ;

  // rule RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_F_T_F_T
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_F_T_F_T =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd5 &&
	     cpReq[61:60] != 2'd2 &&
	     cpReq[9:6] == 4'h9 &&
	     !cpReq[37] &&
	     cpReq_363_BIT_36_924_AND_NOT_wci_busy_5_36_221_ETC___d3245 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_T_T
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_T_T =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     _theResult_____1__h76814 == 4'd5 &&
	     cpReq[37:36] == 2'd2 &&
	     wci_wReset_n_5_16_AND_NOT_wci_busy_5_36_221_AN_ETC___d3224 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_F_T_T
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_F_T_T =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     _theResult_____1__h76814 == 4'd5 &&
	     cpReq[37:36] == 2'd1 &&
	     cpReq[19:9] == 11'd0 &&
	     wci_wReset_n_5_16_AND_NOT_wci_busy_5_36_221_AN_ETC___d3224 ;

  // rule RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_F_T_T_F
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_F_T_T_F =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd6 &&
	     cpReq[61:60] != 2'd2 &&
	     cpReq[9:6] == 4'h9 &&
	     cpReq[37] &&
	     NOT_cpReq_363_BIT_36_924_932_AND_NOT_wci_busy__ETC___d3315 ;

  // rule RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_F_T_F_F
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_F_T_F_F =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd6 &&
	     cpReq[61:60] != 2'd2 &&
	     cpReq[9:6] == 4'h9 &&
	     !cpReq[37] &&
	     NOT_cpReq_363_BIT_36_924_932_AND_NOT_wci_busy__ETC___d3315 ;

  // rule RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_T_T
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_T_T =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd6 &&
	     cpReq[61:60] == 2'd2 &&
	     wci_wReset_n_6_056_AND_NOT_wci_busy_6_076_284__ETC___d3287 ;

  // rule RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_F_T_T_T
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_F_T_T_T =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd6 &&
	     cpReq[61:60] != 2'd2 &&
	     cpReq[9:6] == 4'h9 &&
	     cpReq[37] &&
	     cpReq_363_BIT_36_924_AND_NOT_wci_busy_6_076_28_ETC___d3308 ;

  // rule RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_F_T_F_T
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_F_T_F_T =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd6 &&
	     cpReq[61:60] != 2'd2 &&
	     cpReq[9:6] == 4'h9 &&
	     !cpReq[37] &&
	     cpReq_363_BIT_36_924_AND_NOT_wci_busy_6_076_28_ETC___d3308 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_T_T
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_T_T =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     _theResult_____1__h76814 == 4'd6 &&
	     cpReq[37:36] == 2'd2 &&
	     wci_wReset_n_6_056_AND_NOT_wci_busy_6_076_284__ETC___d3287 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_F_T_T
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_F_T_T =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     _theResult_____1__h76814 == 4'd6 &&
	     cpReq[37:36] == 2'd1 &&
	     cpReq[19:9] == 11'd0 &&
	     wci_wReset_n_6_056_AND_NOT_wci_busy_6_076_284__ETC___d3287 ;

  // rule RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_F_T_T_F
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_F_T_T_F =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd7 &&
	     cpReq[61:60] != 2'd2 &&
	     cpReq[9:6] == 4'h9 &&
	     cpReq[37] &&
	     NOT_cpReq_363_BIT_36_924_932_AND_NOT_wci_busy__ETC___d3378 ;

  // rule RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_F_T_F_F
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_F_T_F_F =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd7 &&
	     cpReq[61:60] != 2'd2 &&
	     cpReq[9:6] == 4'h9 &&
	     !cpReq[37] &&
	     NOT_cpReq_363_BIT_36_924_932_AND_NOT_wci_busy__ETC___d3378 ;

  // rule RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_T_T
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_T_T =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd7 &&
	     cpReq[61:60] == 2'd2 &&
	     wci_wReset_n_7_196_AND_NOT_wci_busy_7_216_347__ETC___d3350 ;

  // rule RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_F_T_T_T
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_F_T_T_T =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd7 &&
	     cpReq[61:60] != 2'd2 &&
	     cpReq[9:6] == 4'h9 &&
	     cpReq[37] &&
	     cpReq_363_BIT_36_924_AND_NOT_wci_busy_7_216_34_ETC___d3371 ;

  // rule RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_F_T_F_T
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_F_T_F_T =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd7 &&
	     cpReq[61:60] != 2'd2 &&
	     cpReq[9:6] == 4'h9 &&
	     !cpReq[37] &&
	     cpReq_363_BIT_36_924_AND_NOT_wci_busy_7_216_34_ETC___d3371 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_T_T
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_T_T =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     _theResult_____1__h76814 == 4'd7 &&
	     cpReq[37:36] == 2'd2 &&
	     wci_wReset_n_7_196_AND_NOT_wci_busy_7_216_347__ETC___d3350 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     _theResult_____1__h76814 == 4'd7 &&
	     cpReq[37:36] == 2'd1 &&
	     cpReq[19:9] == 11'd0 &&
	     wci_wReset_n_7_196_AND_NOT_wci_busy_7_216_347__ETC___d3350 ;

  // rule RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_F_T_T_F
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_F_T_T_F =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd8 &&
	     cpReq[61:60] != 2'd2 &&
	     cpReq[9:6] == 4'h9 &&
	     cpReq[37] &&
	     NOT_cpReq_363_BIT_36_924_932_AND_NOT_wci_busy__ETC___d3441 ;

  // rule RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_F_T_F_F
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_F_T_F_F =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd8 &&
	     cpReq[61:60] != 2'd2 &&
	     cpReq[9:6] == 4'h9 &&
	     !cpReq[37] &&
	     NOT_cpReq_363_BIT_36_924_932_AND_NOT_wci_busy__ETC___d3441 ;

  // rule RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_T_T
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_T_T =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd8 &&
	     cpReq[61:60] == 2'd2 &&
	     wci_wReset_n_8_336_AND_NOT_wci_busy_8_356_410__ETC___d3413 ;

  // rule RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_F_T_T_T
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_F_T_T_T =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd8 &&
	     cpReq[61:60] != 2'd2 &&
	     cpReq[9:6] == 4'h9 &&
	     cpReq[37] &&
	     cpReq_363_BIT_36_924_AND_NOT_wci_busy_8_356_41_ETC___d3434 ;

  // rule RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_F_T_F_T
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_F_T_F_T =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd8 &&
	     cpReq[61:60] != 2'd2 &&
	     cpReq[9:6] == 4'h9 &&
	     !cpReq[37] &&
	     cpReq_363_BIT_36_924_AND_NOT_wci_busy_8_356_41_ETC___d3434 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     _theResult_____1__h76814 == 4'd8 &&
	     cpReq[37:36] == 2'd2 &&
	     wci_wReset_n_8_336_AND_NOT_wci_busy_8_356_410__ETC___d3413 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     _theResult_____1__h76814 == 4'd8 &&
	     cpReq[37:36] == 2'd1 &&
	     cpReq[19:9] == 11'd0 &&
	     wci_wReset_n_8_336_AND_NOT_wci_busy_8_356_410__ETC___d3413 ;

  // rule RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_F_T_T_F
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_F_T_T_F =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd9 &&
	     cpReq[61:60] != 2'd2 &&
	     cpReq[9:6] == 4'h9 &&
	     cpReq[37] &&
	     NOT_cpReq_363_BIT_36_924_932_AND_NOT_wci_busy__ETC___d3504 ;

  // rule RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_F_T_F_F
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_F_T_F_F =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd9 &&
	     cpReq[61:60] != 2'd2 &&
	     cpReq[9:6] == 4'h9 &&
	     !cpReq[37] &&
	     NOT_cpReq_363_BIT_36_924_932_AND_NOT_wci_busy__ETC___d3504 ;

  // rule RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_T_T
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_T_T =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd9 &&
	     cpReq[61:60] == 2'd2 &&
	     wci_wReset_n_9_476_AND_NOT_wci_busy_9_496_473__ETC___d3476 ;

  // rule RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd9 &&
	     cpReq[61:60] != 2'd2 &&
	     cpReq[9:6] == 4'h9 &&
	     cpReq[37] &&
	     cpReq_363_BIT_36_924_AND_NOT_wci_busy_9_496_47_ETC___d3497 ;

  // rule RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_F_T_F_T
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_F_T_F_T =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd9 &&
	     cpReq[61:60] != 2'd2 &&
	     cpReq[9:6] == 4'h9 &&
	     !cpReq[37] &&
	     cpReq_363_BIT_36_924_AND_NOT_wci_busy_9_496_47_ETC___d3497 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     _theResult_____1__h76814 == 4'd9 &&
	     cpReq[37:36] == 2'd2 &&
	     wci_wReset_n_9_476_AND_NOT_wci_busy_9_496_473__ETC___d3476 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     _theResult_____1__h76814 == 4'd9 &&
	     cpReq[37:36] == 2'd1 &&
	     cpReq[19:9] == 11'd0 &&
	     wci_wReset_n_9_476_AND_NOT_wci_busy_9_496_473__ETC___d3476 ;

  // rule RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_F
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_F =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd10 &&
	     cpReq[61:60] != 2'd2 &&
	     cpReq[9:6] == 4'h9 &&
	     cpReq[37] &&
	     NOT_cpReq_363_BIT_36_924_932_AND_NOT_wci_busy__ETC___d3567 ;

  // rule RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_F
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_F =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd10 &&
	     cpReq[61:60] != 2'd2 &&
	     cpReq[9:6] == 4'h9 &&
	     !cpReq[37] &&
	     NOT_cpReq_363_BIT_36_924_932_AND_NOT_wci_busy__ETC___d3567 ;

  // rule RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_T_T
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_T_T =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd10 &&
	     cpReq[61:60] == 2'd2 &&
	     wci_wReset_n_10_616_AND_NOT_wci_busy_10_636_53_ETC___d3539 ;

  // rule RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd10 &&
	     cpReq[61:60] != 2'd2 &&
	     cpReq[9:6] == 4'h9 &&
	     cpReq[37] &&
	     cpReq_363_BIT_36_924_AND_NOT_wci_busy_10_636_5_ETC___d3560 ;

  // rule RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_T
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_T =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd10 &&
	     cpReq[61:60] != 2'd2 &&
	     cpReq[9:6] == 4'h9 &&
	     !cpReq[37] &&
	     cpReq_363_BIT_36_924_AND_NOT_wci_busy_10_636_5_ETC___d3560 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     _theResult_____1__h76814 == 4'd10 &&
	     cpReq[37:36] == 2'd2 &&
	     wci_wReset_n_10_616_AND_NOT_wci_busy_10_636_53_ETC___d3539 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     _theResult_____1__h76814 == 4'd10 &&
	     cpReq[37:36] == 2'd1 &&
	     cpReq[19:9] == 11'd0 &&
	     wci_wReset_n_10_616_AND_NOT_wci_busy_10_636_53_ETC___d3539 ;

  // rule RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_F
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_F =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd11 &&
	     cpReq[61:60] != 2'd2 &&
	     cpReq[9:6] == 4'h9 &&
	     cpReq[37] &&
	     NOT_cpReq_363_BIT_36_924_932_AND_NOT_wci_busy__ETC___d3630 ;

  // rule RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_F
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_F =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd11 &&
	     cpReq[61:60] != 2'd2 &&
	     cpReq[9:6] == 4'h9 &&
	     !cpReq[37] &&
	     NOT_cpReq_363_BIT_36_924_932_AND_NOT_wci_busy__ETC___d3630 ;

  // rule RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_T_T
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_T_T =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd11 &&
	     cpReq[61:60] == 2'd2 &&
	     wci_wReset_n_11_756_AND_NOT_wci_busy_11_776_59_ETC___d3602 ;

  // rule RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd11 &&
	     cpReq[61:60] != 2'd2 &&
	     cpReq[9:6] == 4'h9 &&
	     cpReq[37] &&
	     cpReq_363_BIT_36_924_AND_NOT_wci_busy_11_776_5_ETC___d3623 ;

  // rule RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_T
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_T =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd11 &&
	     cpReq[61:60] != 2'd2 &&
	     cpReq[9:6] == 4'h9 &&
	     !cpReq[37] &&
	     cpReq_363_BIT_36_924_AND_NOT_wci_busy_11_776_5_ETC___d3623 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     _theResult_____1__h76814 == 4'd11 &&
	     cpReq[37:36] == 2'd2 &&
	     wci_wReset_n_11_756_AND_NOT_wci_busy_11_776_59_ETC___d3602 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     _theResult_____1__h76814 == 4'd11 &&
	     cpReq[37:36] == 2'd1 &&
	     cpReq[19:9] == 11'd0 &&
	     wci_wReset_n_11_756_AND_NOT_wci_busy_11_776_59_ETC___d3602 ;

  // rule RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_F
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_F =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd12 &&
	     cpReq[61:60] != 2'd2 &&
	     cpReq[9:6] == 4'h9 &&
	     cpReq[37] &&
	     NOT_cpReq_363_BIT_36_924_932_AND_NOT_wci_busy__ETC___d3693 ;

  // rule RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_F
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_F =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd12 &&
	     cpReq[61:60] != 2'd2 &&
	     cpReq[9:6] == 4'h9 &&
	     !cpReq[37] &&
	     NOT_cpReq_363_BIT_36_924_932_AND_NOT_wci_busy__ETC___d3693 ;

  // rule RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd12 &&
	     cpReq[61:60] == 2'd2 &&
	     wci_wReset_n_12_896_AND_NOT_wci_busy_12_916_66_ETC___d3665 ;

  // rule RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd12 &&
	     cpReq[61:60] != 2'd2 &&
	     cpReq[9:6] == 4'h9 &&
	     cpReq[37] &&
	     cpReq_363_BIT_36_924_AND_NOT_wci_busy_12_916_6_ETC___d3686 ;

  // rule RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_T
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_T =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd12 &&
	     cpReq[61:60] != 2'd2 &&
	     cpReq[9:6] == 4'h9 &&
	     !cpReq[37] &&
	     cpReq_363_BIT_36_924_AND_NOT_wci_busy_12_916_6_ETC___d3686 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     _theResult_____1__h76814 == 4'd12 &&
	     cpReq[37:36] == 2'd2 &&
	     wci_wReset_n_12_896_AND_NOT_wci_busy_12_916_66_ETC___d3665 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     _theResult_____1__h76814 == 4'd12 &&
	     cpReq[37:36] == 2'd1 &&
	     cpReq[19:9] == 11'd0 &&
	     wci_wReset_n_12_896_AND_NOT_wci_busy_12_916_66_ETC___d3665 ;

  // rule RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_F
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_F =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd13 &&
	     cpReq[61:60] != 2'd2 &&
	     cpReq[9:6] == 4'h9 &&
	     cpReq[37] &&
	     NOT_cpReq_363_BIT_36_924_932_AND_NOT_wci_busy__ETC___d3756 ;

  // rule RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_F
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_F =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd13 &&
	     cpReq[61:60] != 2'd2 &&
	     cpReq[9:6] == 4'h9 &&
	     !cpReq[37] &&
	     NOT_cpReq_363_BIT_36_924_932_AND_NOT_wci_busy__ETC___d3756 ;

  // rule RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd13 &&
	     cpReq[61:60] == 2'd2 &&
	     wci_wReset_n_13_036_AND_NOT_wci_busy_13_056_72_ETC___d3728 ;

  // rule RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd13 &&
	     cpReq[61:60] != 2'd2 &&
	     cpReq[9:6] == 4'h9 &&
	     cpReq[37] &&
	     cpReq_363_BIT_36_924_AND_NOT_wci_busy_13_056_7_ETC___d3749 ;

  // rule RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_T
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_T =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd13 &&
	     cpReq[61:60] != 2'd2 &&
	     cpReq[9:6] == 4'h9 &&
	     !cpReq[37] &&
	     cpReq_363_BIT_36_924_AND_NOT_wci_busy_13_056_7_ETC___d3749 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     _theResult_____1__h76814 == 4'd13 &&
	     cpReq[37:36] == 2'd2 &&
	     wci_wReset_n_13_036_AND_NOT_wci_busy_13_056_72_ETC___d3728 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     _theResult_____1__h76814 == 4'd13 &&
	     cpReq[37:36] == 2'd1 &&
	     cpReq[19:9] == 11'd0 &&
	     wci_wReset_n_13_036_AND_NOT_wci_busy_13_056_72_ETC___d3728 ;

  // rule RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_F
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_F =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd14 &&
	     cpReq[61:60] != 2'd2 &&
	     cpReq[9:6] == 4'h9 &&
	     cpReq[37] &&
	     NOT_cpReq_363_BIT_36_924_932_AND_NOT_wci_busy__ETC___d3819 ;

  // rule RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_F
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_F =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd14 &&
	     cpReq[61:60] != 2'd2 &&
	     cpReq[9:6] == 4'h9 &&
	     !cpReq[37] &&
	     NOT_cpReq_363_BIT_36_924_932_AND_NOT_wci_busy__ETC___d3819 ;

  // rule RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd14 &&
	     cpReq[61:60] == 2'd2 &&
	     wci_wReset_n_14_176_AND_NOT_wci_busy_14_196_78_ETC___d3791 ;

  // rule RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd14 &&
	     cpReq[61:60] != 2'd2 &&
	     cpReq[9:6] == 4'h9 &&
	     cpReq[37] &&
	     cpReq_363_BIT_36_924_AND_NOT_wci_busy_14_196_7_ETC___d3812 ;

  // rule RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_T
  assign WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_T =
	     cpReq[64:62] == 3'd3 && _theResult_____1__h76796 == 4'd14 &&
	     cpReq[61:60] != 2'd2 &&
	     cpReq[9:6] == 4'h9 &&
	     !cpReq[37] &&
	     cpReq_363_BIT_36_924_AND_NOT_wci_busy_14_196_7_ETC___d3812 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     _theResult_____1__h76814 == 4'd14 &&
	     cpReq[37:36] == 2'd2 &&
	     wci_wReset_n_14_176_AND_NOT_wci_busy_14_196_78_ETC___d3791 ;

  // rule RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T
  assign WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T =
	     cpReq[64:62] != 3'd1 && cpReq[64:62] != 3'd2 &&
	     cpReq[64:62] != 3'd3 &&
	     cpReq[64:62] != 3'd0 &&
	     _theResult_____1__h76814 == 4'd14 &&
	     cpReq[37:36] == 2'd1 &&
	     cpReq[19:9] == 11'd0 &&
	     wci_wReset_n_14_176_AND_NOT_wci_busy_14_196_78_ETC___d3791 ;

  // rule RL_responseAdminRd
  assign WILL_FIRE_RL_responseAdminRd = adminRespF$EMPTY_N && cpRespF$FULL_N ;

  // rule RL_wci_wrkBusy
  assign WILL_FIRE_RL_wci_wrkBusy =
	     ((wci_wciResponse$wget[33:32] == 2'd0) ?
		wci_respTimr_28_ULT_1_SL_wci_wTimeout_29_30___d5879 ||
		wci_respF$FULL_N :
		wci_respF$FULL_N) &&
	     wci_busy ;

  // rule RL_wci_reqF_incCtr
  assign WILL_FIRE_RL_wci_reqF_incCtr =
	     (wci_reqF_c_r || wci_reqF_x_wire$whas) &&
	     MUX_wci_busy$write_1__SEL_2 &&
	     !wci_reqF_dequeueing$whas ;

  // rule RL_wci_reqF_decCtr
  assign WILL_FIRE_RL_wci_reqF_decCtr =
	     wci_reqF_dequeueing$whas && !MUX_wci_busy$write_1__SEL_2 ;

  // rule RL_wci_reqF_both
  assign WILL_FIRE_RL_wci_reqF_both =
	     (!wci_reqF_c_r || wci_reqF_x_wire$whas) &&
	     wci_reqF_dequeueing$whas &&
	     MUX_wci_busy$write_1__SEL_2 ;

  // rule RL_wci_wrkBusy_1
  assign WILL_FIRE_RL_wci_wrkBusy_1 =
	     ((wci_wciResponse_1$wget[33:32] == 2'd0) ?
		wci_respTimr_1_68_ULT_1_SL_wci_wTimeout_1_69_70___d5880 ||
		wci_respF_1$FULL_N :
		wci_respF_1$FULL_N) &&
	     wci_busy_1 ;

  // rule RL_wci_reqF_1_incCtr
  assign WILL_FIRE_RL_wci_reqF_1_incCtr =
	     (wci_reqF_1_c_r || wci_reqF_1_x_wire$whas) &&
	     MUX_wci_busy_1$write_1__SEL_2 &&
	     !wci_reqF_1_dequeueing$whas ;

  // rule RL_wci_reqF_1_decCtr
  assign WILL_FIRE_RL_wci_reqF_1_decCtr =
	     wci_reqF_1_dequeueing$whas && !MUX_wci_busy_1$write_1__SEL_2 ;

  // rule RL_wci_reqF_1_both
  assign WILL_FIRE_RL_wci_reqF_1_both =
	     (!wci_reqF_1_c_r || wci_reqF_1_x_wire$whas) &&
	     wci_reqF_1_dequeueing$whas &&
	     MUX_wci_busy_1$write_1__SEL_2 ;

  // rule RL_wci_wrkBusy_2
  assign WILL_FIRE_RL_wci_wrkBusy_2 =
	     ((wci_wciResponse_2$wget[33:32] == 2'd0) ?
		wci_respTimr_2_08_ULT_1_SL_wci_wTimeout_2_09_10___d5881 ||
		wci_respF_2$FULL_N :
		wci_respF_2$FULL_N) &&
	     wci_busy_2 ;

  // rule RL_wci_reqF_2_incCtr
  assign WILL_FIRE_RL_wci_reqF_2_incCtr =
	     (wci_reqF_2_c_r || wci_reqF_2_x_wire$whas) &&
	     MUX_wci_busy_2$write_1__SEL_2 &&
	     !wci_reqF_2_dequeueing$whas ;

  // rule RL_wci_reqF_2_decCtr
  assign WILL_FIRE_RL_wci_reqF_2_decCtr =
	     wci_reqF_2_dequeueing$whas && !MUX_wci_busy_2$write_1__SEL_2 ;

  // rule RL_wci_reqF_2_both
  assign WILL_FIRE_RL_wci_reqF_2_both =
	     (!wci_reqF_2_c_r || wci_reqF_2_x_wire$whas) &&
	     wci_reqF_2_dequeueing$whas &&
	     MUX_wci_busy_2$write_1__SEL_2 ;

  // rule RL_wci_wrkBusy_3
  assign WILL_FIRE_RL_wci_wrkBusy_3 =
	     ((wci_wciResponse_3$wget[33:32] == 2'd0) ?
		wci_respTimr_3_48_ULT_1_SL_wci_wTimeout_3_49_50___d5882 ||
		wci_respF_3$FULL_N :
		wci_respF_3$FULL_N) &&
	     wci_busy_3 ;

  // rule RL_wci_reqF_3_incCtr
  assign WILL_FIRE_RL_wci_reqF_3_incCtr =
	     (wci_reqF_3_c_r || wci_reqF_3_x_wire$whas) &&
	     MUX_wci_busy_3$write_1__SEL_2 &&
	     !wci_reqF_3_dequeueing$whas ;

  // rule RL_wci_reqF_3_decCtr
  assign WILL_FIRE_RL_wci_reqF_3_decCtr =
	     wci_reqF_3_dequeueing$whas && !MUX_wci_busy_3$write_1__SEL_2 ;

  // rule RL_wci_reqF_3_both
  assign WILL_FIRE_RL_wci_reqF_3_both =
	     (!wci_reqF_3_c_r || wci_reqF_3_x_wire$whas) &&
	     wci_reqF_3_dequeueing$whas &&
	     MUX_wci_busy_3$write_1__SEL_2 ;

  // rule RL_wci_wrkBusy_4
  assign WILL_FIRE_RL_wci_wrkBusy_4 =
	     ((wci_wciResponse_4$wget[33:32] == 2'd0) ?
		wci_respTimr_4_88_ULT_1_SL_wci_wTimeout_4_89_90___d5883 ||
		wci_respF_4$FULL_N :
		wci_respF_4$FULL_N) &&
	     wci_busy_4 ;

  // rule RL_wci_reqF_4_incCtr
  assign WILL_FIRE_RL_wci_reqF_4_incCtr =
	     (wci_reqF_4_c_r || wci_reqF_4_x_wire$whas) &&
	     MUX_wci_busy_4$write_1__SEL_2 &&
	     !wci_reqF_4_dequeueing$whas ;

  // rule RL_wci_reqF_4_decCtr
  assign WILL_FIRE_RL_wci_reqF_4_decCtr =
	     wci_reqF_4_dequeueing$whas && !MUX_wci_busy_4$write_1__SEL_2 ;

  // rule RL_wci_reqF_4_both
  assign WILL_FIRE_RL_wci_reqF_4_both =
	     (!wci_reqF_4_c_r || wci_reqF_4_x_wire$whas) &&
	     wci_reqF_4_dequeueing$whas &&
	     MUX_wci_busy_4$write_1__SEL_2 ;

  // rule RL_wci_wrkBusy_5
  assign WILL_FIRE_RL_wci_wrkBusy_5 =
	     ((wci_wciResponse_5$wget[33:32] == 2'd0) ?
		wci_respTimr_5_28_ULT_1_SL_wci_wTimeout_5_29_30___d5884 ||
		wci_respF_5$FULL_N :
		wci_respF_5$FULL_N) &&
	     wci_busy_5 ;

  // rule RL_wci_reqF_5_incCtr
  assign WILL_FIRE_RL_wci_reqF_5_incCtr =
	     (wci_reqF_5_c_r || wci_reqF_5_x_wire$whas) &&
	     MUX_wci_busy_5$write_1__SEL_2 &&
	     !wci_reqF_5_dequeueing$whas ;

  // rule RL_wci_reqF_5_decCtr
  assign WILL_FIRE_RL_wci_reqF_5_decCtr =
	     wci_reqF_5_dequeueing$whas && !MUX_wci_busy_5$write_1__SEL_2 ;

  // rule RL_wci_reqF_5_both
  assign WILL_FIRE_RL_wci_reqF_5_both =
	     (!wci_reqF_5_c_r || wci_reqF_5_x_wire$whas) &&
	     wci_reqF_5_dequeueing$whas &&
	     MUX_wci_busy_5$write_1__SEL_2 ;

  // rule RL_wci_wrkBusy_6
  assign WILL_FIRE_RL_wci_wrkBusy_6 =
	     ((wci_wciResponse_6$wget[33:32] == 2'd0) ?
		wci_respTimr_6_068_ULT_1_SL_wci_wTimeout_6_069_ETC___d5885 ||
		wci_respF_6$FULL_N :
		wci_respF_6$FULL_N) &&
	     wci_busy_6 ;

  // rule RL_wci_reqF_6_incCtr
  assign WILL_FIRE_RL_wci_reqF_6_incCtr =
	     (wci_reqF_6_c_r || wci_reqF_6_x_wire$whas) &&
	     MUX_wci_busy_6$write_1__SEL_2 &&
	     !wci_reqF_6_dequeueing$whas ;

  // rule RL_wci_reqF_6_decCtr
  assign WILL_FIRE_RL_wci_reqF_6_decCtr =
	     wci_reqF_6_dequeueing$whas && !MUX_wci_busy_6$write_1__SEL_2 ;

  // rule RL_wci_reqF_6_both
  assign WILL_FIRE_RL_wci_reqF_6_both =
	     (!wci_reqF_6_c_r || wci_reqF_6_x_wire$whas) &&
	     wci_reqF_6_dequeueing$whas &&
	     MUX_wci_busy_6$write_1__SEL_2 ;

  // rule RL_wci_wrkBusy_7
  assign WILL_FIRE_RL_wci_wrkBusy_7 =
	     ((wci_wciResponse_7$wget[33:32] == 2'd0) ?
		wci_respTimr_7_208_ULT_1_SL_wci_wTimeout_7_209_ETC___d5886 ||
		wci_respF_7$FULL_N :
		wci_respF_7$FULL_N) &&
	     wci_busy_7 ;

  // rule RL_wci_reqF_7_incCtr
  assign WILL_FIRE_RL_wci_reqF_7_incCtr =
	     (wci_reqF_7_c_r || wci_reqF_7_x_wire$whas) &&
	     MUX_wci_busy_7$write_1__SEL_2 &&
	     !wci_reqF_7_dequeueing$whas ;

  // rule RL_wci_reqF_7_decCtr
  assign WILL_FIRE_RL_wci_reqF_7_decCtr =
	     wci_reqF_7_dequeueing$whas && !MUX_wci_busy_7$write_1__SEL_2 ;

  // rule RL_wci_reqF_7_both
  assign WILL_FIRE_RL_wci_reqF_7_both =
	     (!wci_reqF_7_c_r || wci_reqF_7_x_wire$whas) &&
	     wci_reqF_7_dequeueing$whas &&
	     MUX_wci_busy_7$write_1__SEL_2 ;

  // rule RL_wci_wrkBusy_8
  assign WILL_FIRE_RL_wci_wrkBusy_8 =
	     ((wci_wciResponse_8$wget[33:32] == 2'd0) ?
		wci_respTimr_8_348_ULT_1_SL_wci_wTimeout_8_349_ETC___d5887 ||
		wci_respF_8$FULL_N :
		wci_respF_8$FULL_N) &&
	     wci_busy_8 ;

  // rule RL_wci_reqF_8_incCtr
  assign WILL_FIRE_RL_wci_reqF_8_incCtr =
	     (wci_reqF_8_c_r || wci_reqF_8_x_wire$whas) &&
	     MUX_wci_busy_8$write_1__SEL_2 &&
	     !wci_reqF_8_dequeueing$whas ;

  // rule RL_wci_reqF_8_decCtr
  assign WILL_FIRE_RL_wci_reqF_8_decCtr =
	     wci_reqF_8_dequeueing$whas && !MUX_wci_busy_8$write_1__SEL_2 ;

  // rule RL_wci_reqF_8_both
  assign WILL_FIRE_RL_wci_reqF_8_both =
	     (!wci_reqF_8_c_r || wci_reqF_8_x_wire$whas) &&
	     wci_reqF_8_dequeueing$whas &&
	     MUX_wci_busy_8$write_1__SEL_2 ;

  // rule RL_wci_wrkBusy_9
  assign WILL_FIRE_RL_wci_wrkBusy_9 =
	     ((wci_wciResponse_9$wget[33:32] == 2'd0) ?
		wci_respTimr_9_488_ULT_1_SL_wci_wTimeout_9_489_ETC___d5888 ||
		wci_respF_9$FULL_N :
		wci_respF_9$FULL_N) &&
	     wci_busy_9 ;

  // rule RL_wci_reqF_9_incCtr
  assign WILL_FIRE_RL_wci_reqF_9_incCtr =
	     (wci_reqF_9_c_r || wci_reqF_9_x_wire$whas) &&
	     MUX_wci_busy_9$write_1__SEL_2 &&
	     !wci_reqF_9_dequeueing$whas ;

  // rule RL_wci_reqF_9_decCtr
  assign WILL_FIRE_RL_wci_reqF_9_decCtr =
	     wci_reqF_9_dequeueing$whas && !MUX_wci_busy_9$write_1__SEL_2 ;

  // rule RL_wci_reqF_9_both
  assign WILL_FIRE_RL_wci_reqF_9_both =
	     (!wci_reqF_9_c_r || wci_reqF_9_x_wire$whas) &&
	     wci_reqF_9_dequeueing$whas &&
	     MUX_wci_busy_9$write_1__SEL_2 ;

  // rule RL_wci_wrkBusy_10
  assign WILL_FIRE_RL_wci_wrkBusy_10 =
	     ((wci_wciResponse_10$wget[33:32] == 2'd0) ?
		wci_respTimr_10_628_ULT_1_SL_wci_wTimeout_10_6_ETC___d5889 ||
		wci_respF_10$FULL_N :
		wci_respF_10$FULL_N) &&
	     wci_busy_10 ;

  // rule RL_wci_reqF_10_incCtr
  assign WILL_FIRE_RL_wci_reqF_10_incCtr =
	     (wci_reqF_10_c_r || wci_reqF_10_x_wire$whas) &&
	     MUX_wci_busy_10$write_1__SEL_2 &&
	     !wci_reqF_10_dequeueing$whas ;

  // rule RL_wci_reqF_10_decCtr
  assign WILL_FIRE_RL_wci_reqF_10_decCtr =
	     wci_reqF_10_dequeueing$whas && !MUX_wci_busy_10$write_1__SEL_2 ;

  // rule RL_wci_reqF_10_both
  assign WILL_FIRE_RL_wci_reqF_10_both =
	     (!wci_reqF_10_c_r || wci_reqF_10_x_wire$whas) &&
	     wci_reqF_10_dequeueing$whas &&
	     MUX_wci_busy_10$write_1__SEL_2 ;

  // rule RL_wci_wrkBusy_11
  assign WILL_FIRE_RL_wci_wrkBusy_11 =
	     ((wci_wciResponse_11$wget[33:32] == 2'd0) ?
		wci_respTimr_11_768_ULT_1_SL_wci_wTimeout_11_7_ETC___d5890 ||
		wci_respF_11$FULL_N :
		wci_respF_11$FULL_N) &&
	     wci_busy_11 ;

  // rule RL_wci_reqF_11_incCtr
  assign WILL_FIRE_RL_wci_reqF_11_incCtr =
	     (wci_reqF_11_c_r || wci_reqF_11_x_wire$whas) &&
	     MUX_wci_busy_11$write_1__SEL_2 &&
	     !wci_reqF_11_dequeueing$whas ;

  // rule RL_wci_reqF_11_decCtr
  assign WILL_FIRE_RL_wci_reqF_11_decCtr =
	     wci_reqF_11_dequeueing$whas && !MUX_wci_busy_11$write_1__SEL_2 ;

  // rule RL_wci_reqF_11_both
  assign WILL_FIRE_RL_wci_reqF_11_both =
	     (!wci_reqF_11_c_r || wci_reqF_11_x_wire$whas) &&
	     wci_reqF_11_dequeueing$whas &&
	     MUX_wci_busy_11$write_1__SEL_2 ;

  // rule RL_wci_wrkBusy_12
  assign WILL_FIRE_RL_wci_wrkBusy_12 =
	     ((wci_wciResponse_12$wget[33:32] == 2'd0) ?
		wci_respTimr_12_908_ULT_1_SL_wci_wTimeout_12_9_ETC___d5891 ||
		wci_respF_12$FULL_N :
		wci_respF_12$FULL_N) &&
	     wci_busy_12 ;

  // rule RL_wci_reqF_12_incCtr
  assign WILL_FIRE_RL_wci_reqF_12_incCtr =
	     (wci_reqF_12_c_r || wci_reqF_12_x_wire$whas) &&
	     MUX_wci_busy_12$write_1__SEL_2 &&
	     !wci_reqF_12_dequeueing$whas ;

  // rule RL_wci_reqF_12_decCtr
  assign WILL_FIRE_RL_wci_reqF_12_decCtr =
	     wci_reqF_12_dequeueing$whas && !MUX_wci_busy_12$write_1__SEL_2 ;

  // rule RL_wci_reqF_12_both
  assign WILL_FIRE_RL_wci_reqF_12_both =
	     (!wci_reqF_12_c_r || wci_reqF_12_x_wire$whas) &&
	     wci_reqF_12_dequeueing$whas &&
	     MUX_wci_busy_12$write_1__SEL_2 ;

  // rule RL_wci_wrkBusy_13
  assign WILL_FIRE_RL_wci_wrkBusy_13 =
	     ((wci_wciResponse_13$wget[33:32] == 2'd0) ?
		wci_respTimr_13_048_ULT_1_SL_wci_wTimeout_13_0_ETC___d5892 ||
		wci_respF_13$FULL_N :
		wci_respF_13$FULL_N) &&
	     wci_busy_13 ;

  // rule RL_wci_reqF_13_incCtr
  assign WILL_FIRE_RL_wci_reqF_13_incCtr =
	     (wci_reqF_13_c_r || wci_reqF_13_x_wire$whas) &&
	     MUX_wci_busy_13$write_1__SEL_2 &&
	     !wci_reqF_13_dequeueing$whas ;

  // rule RL_wci_reqF_13_decCtr
  assign WILL_FIRE_RL_wci_reqF_13_decCtr =
	     wci_reqF_13_dequeueing$whas && !MUX_wci_busy_13$write_1__SEL_2 ;

  // rule RL_wci_reqF_13_both
  assign WILL_FIRE_RL_wci_reqF_13_both =
	     (!wci_reqF_13_c_r || wci_reqF_13_x_wire$whas) &&
	     wci_reqF_13_dequeueing$whas &&
	     MUX_wci_busy_13$write_1__SEL_2 ;

  // rule RL_wci_wrkBusy_14
  assign WILL_FIRE_RL_wci_wrkBusy_14 =
	     ((wci_wciResponse_14$wget[33:32] == 2'd0) ?
		wci_respTimr_14_188_ULT_1_SL_wci_wTimeout_14_1_ETC___d5893 ||
		wci_respF_14$FULL_N :
		wci_respF_14$FULL_N) &&
	     wci_busy_14 ;

  // rule RL_wci_reqF_14_incCtr
  assign WILL_FIRE_RL_wci_reqF_14_incCtr =
	     (wci_reqF_14_c_r || wci_reqF_14_x_wire$whas) &&
	     MUX_wci_busy_14$write_1__SEL_2 &&
	     !wci_reqF_14_dequeueing$whas ;

  // rule RL_wci_reqF_14_decCtr
  assign WILL_FIRE_RL_wci_reqF_14_decCtr =
	     wci_reqF_14_dequeueing$whas && !MUX_wci_busy_14$write_1__SEL_2 ;

  // rule RL_wci_reqF_14_both
  assign WILL_FIRE_RL_wci_reqF_14_both =
	     (!wci_reqF_14_c_r || wci_reqF_14_x_wire$whas) &&
	     wci_reqF_14_dequeueing$whas &&
	     MUX_wci_busy_14$write_1__SEL_2 ;

  // inputs to muxes for submodule ports
  assign MUX_wci_busy$write_1__SEL_1 =
	     WILL_FIRE_RL_wci_wrkBusy &&
	     (!wci_respTimr_28_ULT_1_SL_wci_wTimeout_29_30___d5879 ||
	      wci_wciResponse$wget[33:32] != 2'd0) ;
  assign MUX_wci_busy$write_1__SEL_2 =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_T_F_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_T_T_T ;
  assign MUX_wci_busy_1$write_1__SEL_1 =
	     WILL_FIRE_RL_wci_wrkBusy_1 &&
	     (!wci_respTimr_1_68_ULT_1_SL_wci_wTimeout_1_69_70___d5880 ||
	      wci_wciResponse_1$wget[33:32] != 2'd0) ;
  assign MUX_wci_busy_1$write_1__SEL_2 =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_F_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_T_T_T ;
  assign MUX_wci_busy_10$write_1__SEL_1 =
	     WILL_FIRE_RL_wci_wrkBusy_10 &&
	     (!wci_respTimr_10_628_ULT_1_SL_wci_wTimeout_10_6_ETC___d5889 ||
	      wci_wciResponse_10$wget[33:32] != 2'd0) ;
  assign MUX_wci_busy_10$write_1__SEL_2 =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_T_T ;
  assign MUX_wci_busy_11$write_1__SEL_1 =
	     WILL_FIRE_RL_wci_wrkBusy_11 &&
	     (!wci_respTimr_11_768_ULT_1_SL_wci_wTimeout_11_7_ETC___d5890 ||
	      wci_wciResponse_11$wget[33:32] != 2'd0) ;
  assign MUX_wci_busy_11$write_1__SEL_2 =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_T_T ;
  assign MUX_wci_busy_12$write_1__SEL_1 =
	     WILL_FIRE_RL_wci_wrkBusy_12 &&
	     (!wci_respTimr_12_908_ULT_1_SL_wci_wTimeout_12_9_ETC___d5891 ||
	      wci_wciResponse_12$wget[33:32] != 2'd0) ;
  assign MUX_wci_busy_12$write_1__SEL_2 =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ;
  assign MUX_wci_busy_13$write_1__SEL_1 =
	     WILL_FIRE_RL_wci_wrkBusy_13 &&
	     (!wci_respTimr_13_048_ULT_1_SL_wci_wTimeout_13_0_ETC___d5892 ||
	      wci_wciResponse_13$wget[33:32] != 2'd0) ;
  assign MUX_wci_busy_13$write_1__SEL_2 =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ;
  assign MUX_wci_busy_14$write_1__SEL_1 =
	     WILL_FIRE_RL_wci_wrkBusy_14 &&
	     (!wci_respTimr_14_188_ULT_1_SL_wci_wTimeout_14_1_ETC___d5893 ||
	      wci_wciResponse_14$wget[33:32] != 2'd0) ;
  assign MUX_wci_busy_14$write_1__SEL_2 =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ;
  assign MUX_wci_busy_2$write_1__SEL_1 =
	     WILL_FIRE_RL_wci_wrkBusy_2 &&
	     (!wci_respTimr_2_08_ULT_1_SL_wci_wTimeout_2_09_10___d5881 ||
	      wci_wciResponse_2$wget[33:32] != 2'd0) ;
  assign MUX_wci_busy_2$write_1__SEL_2 =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_F_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_T_T ;
  assign MUX_wci_busy_3$write_1__SEL_1 =
	     WILL_FIRE_RL_wci_wrkBusy_3 &&
	     (!wci_respTimr_3_48_ULT_1_SL_wci_wTimeout_3_49_50___d5882 ||
	      wci_wciResponse_3$wget[33:32] != 2'd0) ;
  assign MUX_wci_busy_3$write_1__SEL_2 =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_F_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_T_T ;
  assign MUX_wci_busy_4$write_1__SEL_1 =
	     WILL_FIRE_RL_wci_wrkBusy_4 &&
	     (!wci_respTimr_4_88_ULT_1_SL_wci_wTimeout_4_89_90___d5883 ||
	      wci_wciResponse_4$wget[33:32] != 2'd0) ;
  assign MUX_wci_busy_4$write_1__SEL_2 =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_F_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_T_T ;
  assign MUX_wci_busy_5$write_1__SEL_1 =
	     WILL_FIRE_RL_wci_wrkBusy_5 &&
	     (!wci_respTimr_5_28_ULT_1_SL_wci_wTimeout_5_29_30___d5884 ||
	      wci_wciResponse_5$wget[33:32] != 2'd0) ;
  assign MUX_wci_busy_5$write_1__SEL_2 =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_F_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_T_T ;
  assign MUX_wci_busy_6$write_1__SEL_1 =
	     WILL_FIRE_RL_wci_wrkBusy_6 &&
	     (!wci_respTimr_6_068_ULT_1_SL_wci_wTimeout_6_069_ETC___d5885 ||
	      wci_wciResponse_6$wget[33:32] != 2'd0) ;
  assign MUX_wci_busy_6$write_1__SEL_2 =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_F_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_T_T ;
  assign MUX_wci_busy_7$write_1__SEL_1 =
	     WILL_FIRE_RL_wci_wrkBusy_7 &&
	     (!wci_respTimr_7_208_ULT_1_SL_wci_wTimeout_7_209_ETC___d5886 ||
	      wci_wciResponse_7$wget[33:32] != 2'd0) ;
  assign MUX_wci_busy_7$write_1__SEL_2 =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_T_T ;
  assign MUX_wci_busy_8$write_1__SEL_1 =
	     WILL_FIRE_RL_wci_wrkBusy_8 &&
	     (!wci_respTimr_8_348_ULT_1_SL_wci_wTimeout_8_349_ETC___d5887 ||
	      wci_wciResponse_8$wget[33:32] != 2'd0) ;
  assign MUX_wci_busy_8$write_1__SEL_2 =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_T_T ;
  assign MUX_wci_busy_9$write_1__SEL_1 =
	     WILL_FIRE_RL_wci_wrkBusy_9 &&
	     (!wci_respTimr_9_488_ULT_1_SL_wci_wTimeout_9_489_ETC___d5888 ||
	      wci_wciResponse_9$wget[33:32] != 2'd0) ;
  assign MUX_wci_busy_9$write_1__SEL_2 =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_T_T ;
  assign MUX_wci_reqERR$write_1__SEL_1 =
	     WILL_FIRE_RL_wci_wrkBusy &&
	     wci_wciResponse$wget[33:32] == 2'd3 &&
	     (wci_reqPend == 2'd1 || wci_reqPend == 2'd2 ||
	      wci_reqPend == 2'd3) ;
  assign MUX_wci_reqERR_1$write_1__SEL_1 =
	     WILL_FIRE_RL_wci_wrkBusy_1 &&
	     wci_wciResponse_1$wget[33:32] == 2'd3 &&
	     (wci_reqPend_1 == 2'd1 || wci_reqPend_1 == 2'd2 ||
	      wci_reqPend_1 == 2'd3) ;
  assign MUX_wci_reqERR_10$write_1__SEL_1 =
	     WILL_FIRE_RL_wci_wrkBusy_10 &&
	     wci_wciResponse_10$wget[33:32] == 2'd3 &&
	     (wci_reqPend_10 == 2'd1 || wci_reqPend_10 == 2'd2 ||
	      wci_reqPend_10 == 2'd3) ;
  assign MUX_wci_reqERR_11$write_1__SEL_1 =
	     WILL_FIRE_RL_wci_wrkBusy_11 &&
	     wci_wciResponse_11$wget[33:32] == 2'd3 &&
	     (wci_reqPend_11 == 2'd1 || wci_reqPend_11 == 2'd2 ||
	      wci_reqPend_11 == 2'd3) ;
  assign MUX_wci_reqERR_12$write_1__SEL_1 =
	     WILL_FIRE_RL_wci_wrkBusy_12 &&
	     wci_wciResponse_12$wget[33:32] == 2'd3 &&
	     (wci_reqPend_12 == 2'd1 || wci_reqPend_12 == 2'd2 ||
	      wci_reqPend_12 == 2'd3) ;
  assign MUX_wci_reqERR_13$write_1__SEL_1 =
	     WILL_FIRE_RL_wci_wrkBusy_13 &&
	     wci_wciResponse_13$wget[33:32] == 2'd3 &&
	     (wci_reqPend_13 == 2'd1 || wci_reqPend_13 == 2'd2 ||
	      wci_reqPend_13 == 2'd3) ;
  assign MUX_wci_reqERR_14$write_1__SEL_1 =
	     WILL_FIRE_RL_wci_wrkBusy_14 &&
	     wci_wciResponse_14$wget[33:32] == 2'd3 &&
	     (wci_reqPend_14 == 2'd1 || wci_reqPend_14 == 2'd2 ||
	      wci_reqPend_14 == 2'd3) ;
  assign MUX_wci_reqERR_2$write_1__SEL_1 =
	     WILL_FIRE_RL_wci_wrkBusy_2 &&
	     wci_wciResponse_2$wget[33:32] == 2'd3 &&
	     (wci_reqPend_2 == 2'd1 || wci_reqPend_2 == 2'd2 ||
	      wci_reqPend_2 == 2'd3) ;
  assign MUX_wci_reqERR_3$write_1__SEL_1 =
	     WILL_FIRE_RL_wci_wrkBusy_3 &&
	     wci_wciResponse_3$wget[33:32] == 2'd3 &&
	     (wci_reqPend_3 == 2'd1 || wci_reqPend_3 == 2'd2 ||
	      wci_reqPend_3 == 2'd3) ;
  assign MUX_wci_reqERR_4$write_1__SEL_1 =
	     WILL_FIRE_RL_wci_wrkBusy_4 &&
	     wci_wciResponse_4$wget[33:32] == 2'd3 &&
	     (wci_reqPend_4 == 2'd1 || wci_reqPend_4 == 2'd2 ||
	      wci_reqPend_4 == 2'd3) ;
  assign MUX_wci_reqERR_5$write_1__SEL_1 =
	     WILL_FIRE_RL_wci_wrkBusy_5 &&
	     wci_wciResponse_5$wget[33:32] == 2'd3 &&
	     (wci_reqPend_5 == 2'd1 || wci_reqPend_5 == 2'd2 ||
	      wci_reqPend_5 == 2'd3) ;
  assign MUX_wci_reqERR_6$write_1__SEL_1 =
	     WILL_FIRE_RL_wci_wrkBusy_6 &&
	     wci_wciResponse_6$wget[33:32] == 2'd3 &&
	     (wci_reqPend_6 == 2'd1 || wci_reqPend_6 == 2'd2 ||
	      wci_reqPend_6 == 2'd3) ;
  assign MUX_wci_reqERR_7$write_1__SEL_1 =
	     WILL_FIRE_RL_wci_wrkBusy_7 &&
	     wci_wciResponse_7$wget[33:32] == 2'd3 &&
	     (wci_reqPend_7 == 2'd1 || wci_reqPend_7 == 2'd2 ||
	      wci_reqPend_7 == 2'd3) ;
  assign MUX_wci_reqERR_8$write_1__SEL_1 =
	     WILL_FIRE_RL_wci_wrkBusy_8 &&
	     wci_wciResponse_8$wget[33:32] == 2'd3 &&
	     (wci_reqPend_8 == 2'd1 || wci_reqPend_8 == 2'd2 ||
	      wci_reqPend_8 == 2'd3) ;
  assign MUX_wci_reqERR_9$write_1__SEL_1 =
	     WILL_FIRE_RL_wci_wrkBusy_9 &&
	     wci_wciResponse_9$wget[33:32] == 2'd3 &&
	     (wci_reqPend_9 == 2'd1 || wci_reqPend_9 == 2'd2 ||
	      wci_reqPend_9 == 2'd3) ;
  assign MUX_wci_reqFAIL$write_1__SEL_1 =
	     WILL_FIRE_RL_wci_wrkBusy &&
	     wci_wciResponse$wget[33:32] == 2'd2 &&
	     (wci_reqPend == 2'd1 || wci_reqPend == 2'd2 ||
	      wci_reqPend == 2'd3) ;
  assign MUX_wci_reqFAIL_1$write_1__SEL_1 =
	     WILL_FIRE_RL_wci_wrkBusy_1 &&
	     wci_wciResponse_1$wget[33:32] == 2'd2 &&
	     (wci_reqPend_1 == 2'd1 || wci_reqPend_1 == 2'd2 ||
	      wci_reqPend_1 == 2'd3) ;
  assign MUX_wci_reqFAIL_10$write_1__SEL_1 =
	     WILL_FIRE_RL_wci_wrkBusy_10 &&
	     wci_wciResponse_10$wget[33:32] == 2'd2 &&
	     (wci_reqPend_10 == 2'd1 || wci_reqPend_10 == 2'd2 ||
	      wci_reqPend_10 == 2'd3) ;
  assign MUX_wci_reqFAIL_11$write_1__SEL_1 =
	     WILL_FIRE_RL_wci_wrkBusy_11 &&
	     wci_wciResponse_11$wget[33:32] == 2'd2 &&
	     (wci_reqPend_11 == 2'd1 || wci_reqPend_11 == 2'd2 ||
	      wci_reqPend_11 == 2'd3) ;
  assign MUX_wci_reqFAIL_12$write_1__SEL_1 =
	     WILL_FIRE_RL_wci_wrkBusy_12 &&
	     wci_wciResponse_12$wget[33:32] == 2'd2 &&
	     (wci_reqPend_12 == 2'd1 || wci_reqPend_12 == 2'd2 ||
	      wci_reqPend_12 == 2'd3) ;
  assign MUX_wci_reqFAIL_13$write_1__SEL_1 =
	     WILL_FIRE_RL_wci_wrkBusy_13 &&
	     wci_wciResponse_13$wget[33:32] == 2'd2 &&
	     (wci_reqPend_13 == 2'd1 || wci_reqPend_13 == 2'd2 ||
	      wci_reqPend_13 == 2'd3) ;
  assign MUX_wci_reqFAIL_14$write_1__SEL_1 =
	     WILL_FIRE_RL_wci_wrkBusy_14 &&
	     wci_wciResponse_14$wget[33:32] == 2'd2 &&
	     (wci_reqPend_14 == 2'd1 || wci_reqPend_14 == 2'd2 ||
	      wci_reqPend_14 == 2'd3) ;
  assign MUX_wci_reqFAIL_2$write_1__SEL_1 =
	     WILL_FIRE_RL_wci_wrkBusy_2 &&
	     wci_wciResponse_2$wget[33:32] == 2'd2 &&
	     (wci_reqPend_2 == 2'd1 || wci_reqPend_2 == 2'd2 ||
	      wci_reqPend_2 == 2'd3) ;
  assign MUX_wci_reqFAIL_3$write_1__SEL_1 =
	     WILL_FIRE_RL_wci_wrkBusy_3 &&
	     wci_wciResponse_3$wget[33:32] == 2'd2 &&
	     (wci_reqPend_3 == 2'd1 || wci_reqPend_3 == 2'd2 ||
	      wci_reqPend_3 == 2'd3) ;
  assign MUX_wci_reqFAIL_4$write_1__SEL_1 =
	     WILL_FIRE_RL_wci_wrkBusy_4 &&
	     wci_wciResponse_4$wget[33:32] == 2'd2 &&
	     (wci_reqPend_4 == 2'd1 || wci_reqPend_4 == 2'd2 ||
	      wci_reqPend_4 == 2'd3) ;
  assign MUX_wci_reqFAIL_5$write_1__SEL_1 =
	     WILL_FIRE_RL_wci_wrkBusy_5 &&
	     wci_wciResponse_5$wget[33:32] == 2'd2 &&
	     (wci_reqPend_5 == 2'd1 || wci_reqPend_5 == 2'd2 ||
	      wci_reqPend_5 == 2'd3) ;
  assign MUX_wci_reqFAIL_6$write_1__SEL_1 =
	     WILL_FIRE_RL_wci_wrkBusy_6 &&
	     wci_wciResponse_6$wget[33:32] == 2'd2 &&
	     (wci_reqPend_6 == 2'd1 || wci_reqPend_6 == 2'd2 ||
	      wci_reqPend_6 == 2'd3) ;
  assign MUX_wci_reqFAIL_7$write_1__SEL_1 =
	     WILL_FIRE_RL_wci_wrkBusy_7 &&
	     wci_wciResponse_7$wget[33:32] == 2'd2 &&
	     (wci_reqPend_7 == 2'd1 || wci_reqPend_7 == 2'd2 ||
	      wci_reqPend_7 == 2'd3) ;
  assign MUX_wci_reqFAIL_8$write_1__SEL_1 =
	     WILL_FIRE_RL_wci_wrkBusy_8 &&
	     wci_wciResponse_8$wget[33:32] == 2'd2 &&
	     (wci_reqPend_8 == 2'd1 || wci_reqPend_8 == 2'd2 ||
	      wci_reqPend_8 == 2'd3) ;
  assign MUX_wci_reqFAIL_9$write_1__SEL_1 =
	     WILL_FIRE_RL_wci_wrkBusy_9 &&
	     wci_wciResponse_9$wget[33:32] == 2'd2 &&
	     (wci_reqPend_9 == 2'd1 || wci_reqPend_9 == 2'd2 ||
	      wci_reqPend_9 == 2'd3) ;
  assign MUX_wci_reqF_10_q_0$write_1__SEL_1 =
	     WILL_FIRE_RL_wci_reqF_10_incCtr && !wci_reqF_10_c_r ;
  assign MUX_wci_reqF_11_q_0$write_1__SEL_1 =
	     WILL_FIRE_RL_wci_reqF_11_incCtr && !wci_reqF_11_c_r ;
  assign MUX_wci_reqF_12_q_0$write_1__SEL_1 =
	     WILL_FIRE_RL_wci_reqF_12_incCtr && !wci_reqF_12_c_r ;
  assign MUX_wci_reqF_13_q_0$write_1__SEL_1 =
	     WILL_FIRE_RL_wci_reqF_13_incCtr && !wci_reqF_13_c_r ;
  assign MUX_wci_reqF_14_q_0$write_1__SEL_1 =
	     WILL_FIRE_RL_wci_reqF_14_incCtr && !wci_reqF_14_c_r ;
  assign MUX_wci_reqF_1_q_0$write_1__SEL_2 =
	     WILL_FIRE_RL_wci_reqF_1_incCtr && !wci_reqF_1_c_r ;
  assign MUX_wci_reqF_2_q_0$write_1__SEL_2 =
	     WILL_FIRE_RL_wci_reqF_2_incCtr && !wci_reqF_2_c_r ;
  assign MUX_wci_reqF_3_q_0$write_1__SEL_2 =
	     WILL_FIRE_RL_wci_reqF_3_incCtr && !wci_reqF_3_c_r ;
  assign MUX_wci_reqF_4_q_0$write_1__SEL_2 =
	     WILL_FIRE_RL_wci_reqF_4_incCtr && !wci_reqF_4_c_r ;
  assign MUX_wci_reqF_5_q_0$write_1__SEL_2 =
	     WILL_FIRE_RL_wci_reqF_5_incCtr && !wci_reqF_5_c_r ;
  assign MUX_wci_reqF_6_q_0$write_1__SEL_2 =
	     WILL_FIRE_RL_wci_reqF_6_incCtr && !wci_reqF_6_c_r ;
  assign MUX_wci_reqF_7_q_0$write_1__SEL_2 =
	     WILL_FIRE_RL_wci_reqF_7_incCtr && !wci_reqF_7_c_r ;
  assign MUX_wci_reqF_8_q_0$write_1__SEL_2 =
	     WILL_FIRE_RL_wci_reqF_8_incCtr && !wci_reqF_8_c_r ;
  assign MUX_wci_reqF_9_q_0$write_1__SEL_2 =
	     WILL_FIRE_RL_wci_reqF_9_incCtr && !wci_reqF_9_c_r ;
  assign MUX_wci_reqF_q_0$write_1__SEL_2 =
	     WILL_FIRE_RL_wci_reqF_incCtr && !wci_reqF_c_r ;
  assign MUX_wci_reqPend$write_1__SEL_1 =
	     WILL_FIRE_RL_wci_wrkBusy && wci_wciResponse$wget[33:32] != 2'd0 ;
  assign MUX_wci_reqPend_1$write_1__SEL_1 =
	     WILL_FIRE_RL_wci_wrkBusy_1 &&
	     wci_wciResponse_1$wget[33:32] != 2'd0 ;
  assign MUX_wci_reqPend_10$write_1__SEL_1 =
	     WILL_FIRE_RL_wci_wrkBusy_10 &&
	     wci_wciResponse_10$wget[33:32] != 2'd0 ;
  assign MUX_wci_reqPend_11$write_1__SEL_1 =
	     WILL_FIRE_RL_wci_wrkBusy_11 &&
	     wci_wciResponse_11$wget[33:32] != 2'd0 ;
  assign MUX_wci_reqPend_12$write_1__SEL_1 =
	     WILL_FIRE_RL_wci_wrkBusy_12 &&
	     wci_wciResponse_12$wget[33:32] != 2'd0 ;
  assign MUX_wci_reqPend_13$write_1__SEL_1 =
	     WILL_FIRE_RL_wci_wrkBusy_13 &&
	     wci_wciResponse_13$wget[33:32] != 2'd0 ;
  assign MUX_wci_reqPend_14$write_1__SEL_1 =
	     WILL_FIRE_RL_wci_wrkBusy_14 &&
	     wci_wciResponse_14$wget[33:32] != 2'd0 ;
  assign MUX_wci_reqPend_2$write_1__SEL_1 =
	     WILL_FIRE_RL_wci_wrkBusy_2 &&
	     wci_wciResponse_2$wget[33:32] != 2'd0 ;
  assign MUX_wci_reqPend_3$write_1__SEL_1 =
	     WILL_FIRE_RL_wci_wrkBusy_3 &&
	     wci_wciResponse_3$wget[33:32] != 2'd0 ;
  assign MUX_wci_reqPend_4$write_1__SEL_1 =
	     WILL_FIRE_RL_wci_wrkBusy_4 &&
	     wci_wciResponse_4$wget[33:32] != 2'd0 ;
  assign MUX_wci_reqPend_5$write_1__SEL_1 =
	     WILL_FIRE_RL_wci_wrkBusy_5 &&
	     wci_wciResponse_5$wget[33:32] != 2'd0 ;
  assign MUX_wci_reqPend_6$write_1__SEL_1 =
	     WILL_FIRE_RL_wci_wrkBusy_6 &&
	     wci_wciResponse_6$wget[33:32] != 2'd0 ;
  assign MUX_wci_reqPend_7$write_1__SEL_1 =
	     WILL_FIRE_RL_wci_wrkBusy_7 &&
	     wci_wciResponse_7$wget[33:32] != 2'd0 ;
  assign MUX_wci_reqPend_8$write_1__SEL_1 =
	     WILL_FIRE_RL_wci_wrkBusy_8 &&
	     wci_wciResponse_8$wget[33:32] != 2'd0 ;
  assign MUX_wci_reqPend_9$write_1__SEL_1 =
	     WILL_FIRE_RL_wci_wrkBusy_9 &&
	     wci_wciResponse_9$wget[33:32] != 2'd0 ;
  assign MUX_wci_reqTO$write_1__SEL_1 =
	     WILL_FIRE_RL_wci_wrkBusy &&
	     wci_wciResponse_wget__23_BITS_33_TO_32_24_EQ_0_ETC___d252 ;
  assign MUX_wci_reqTO_1$write_1__SEL_1 =
	     WILL_FIRE_RL_wci_wrkBusy_1 &&
	     wci_wciResponse_1_wget__63_BITS_33_TO_32_64_EQ_ETC___d392 ;
  assign MUX_wci_reqTO_10$write_1__SEL_1 =
	     WILL_FIRE_RL_wci_wrkBusy_10 &&
	     wci_wciResponse_10_wget__623_BITS_33_TO_32_624_ETC___d1652 ;
  assign MUX_wci_reqTO_11$write_1__SEL_1 =
	     WILL_FIRE_RL_wci_wrkBusy_11 &&
	     wci_wciResponse_11_wget__763_BITS_33_TO_32_764_ETC___d1792 ;
  assign MUX_wci_reqTO_12$write_1__SEL_1 =
	     WILL_FIRE_RL_wci_wrkBusy_12 &&
	     wci_wciResponse_12_wget__903_BITS_33_TO_32_904_ETC___d1932 ;
  assign MUX_wci_reqTO_13$write_1__SEL_1 =
	     WILL_FIRE_RL_wci_wrkBusy_13 &&
	     wci_wciResponse_13_wget__043_BITS_33_TO_32_044_ETC___d2072 ;
  assign MUX_wci_reqTO_14$write_1__SEL_1 =
	     WILL_FIRE_RL_wci_wrkBusy_14 &&
	     wci_wciResponse_14_wget__183_BITS_33_TO_32_184_ETC___d2212 ;
  assign MUX_wci_reqTO_2$write_1__SEL_1 =
	     WILL_FIRE_RL_wci_wrkBusy_2 &&
	     wci_wciResponse_2_wget__03_BITS_33_TO_32_04_EQ_ETC___d532 ;
  assign MUX_wci_reqTO_3$write_1__SEL_1 =
	     WILL_FIRE_RL_wci_wrkBusy_3 &&
	     wci_wciResponse_3_wget__43_BITS_33_TO_32_44_EQ_ETC___d672 ;
  assign MUX_wci_reqTO_4$write_1__SEL_1 =
	     WILL_FIRE_RL_wci_wrkBusy_4 &&
	     wci_wciResponse_4_wget__83_BITS_33_TO_32_84_EQ_ETC___d812 ;
  assign MUX_wci_reqTO_5$write_1__SEL_1 =
	     WILL_FIRE_RL_wci_wrkBusy_5 &&
	     wci_wciResponse_5_wget__23_BITS_33_TO_32_24_EQ_ETC___d952 ;
  assign MUX_wci_reqTO_6$write_1__SEL_1 =
	     WILL_FIRE_RL_wci_wrkBusy_6 &&
	     wci_wciResponse_6_wget__063_BITS_33_TO_32_064__ETC___d1092 ;
  assign MUX_wci_reqTO_7$write_1__SEL_1 =
	     WILL_FIRE_RL_wci_wrkBusy_7 &&
	     wci_wciResponse_7_wget__203_BITS_33_TO_32_204__ETC___d1232 ;
  assign MUX_wci_reqTO_8$write_1__SEL_1 =
	     WILL_FIRE_RL_wci_wrkBusy_8 &&
	     wci_wciResponse_8_wget__343_BITS_33_TO_32_344__ETC___d1372 ;
  assign MUX_wci_reqTO_9$write_1__SEL_1 =
	     WILL_FIRE_RL_wci_wrkBusy_9 &&
	     wci_wciResponse_9_wget__483_BITS_33_TO_32_484__ETC___d1512 ;
  assign MUX_wci_respF$enq_1__SEL_6 =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_T_F_F_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_T_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_T_F_F_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_T_F_F_T_T_T ;
  assign MUX_wci_respF$enq_1__SEL_7 =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_T_F_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_T_T_F ;
  assign MUX_wci_respF_1$enq_1__SEL_6 =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_F_F_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_T_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_T_F_F_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_T_F_F_T_T_T ;
  assign MUX_wci_respF_1$enq_1__SEL_7 =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_F_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_T_T_F ;
  assign MUX_wci_respF_10$enq_1__SEL_6 =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T ;
  assign MUX_wci_respF_10$enq_1__SEL_7 =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_T_F ;
  assign MUX_wci_respF_11$enq_1__SEL_6 =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T ;
  assign MUX_wci_respF_11$enq_1__SEL_7 =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_T_F ;
  assign MUX_wci_respF_12$enq_1__SEL_6 =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T ;
  assign MUX_wci_respF_12$enq_1__SEL_7 =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F ;
  assign MUX_wci_respF_13$enq_1__SEL_6 =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T ;
  assign MUX_wci_respF_13$enq_1__SEL_7 =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F ;
  assign MUX_wci_respF_14$enq_1__SEL_6 =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T ;
  assign MUX_wci_respF_14$enq_1__SEL_7 =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F ;
  assign MUX_wci_respF_2$enq_1__SEL_6 =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_F_F_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_F_F_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_F_F_T_T_T ;
  assign MUX_wci_respF_2$enq_1__SEL_7 =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_F_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_T_F ;
  assign MUX_wci_respF_3$enq_1__SEL_6 =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_F_F_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_F_F_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_F_F_T_T_T ;
  assign MUX_wci_respF_3$enq_1__SEL_7 =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_F_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_T_F ;
  assign MUX_wci_respF_4$enq_1__SEL_6 =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_F_F_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_F_F_T_T_T ;
  assign MUX_wci_respF_4$enq_1__SEL_7 =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_F_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_T_F ;
  assign MUX_wci_respF_5$enq_1__SEL_6 =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_F_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_F_T_T_T ;
  assign MUX_wci_respF_5$enq_1__SEL_7 =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_F_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_T_F ;
  assign MUX_wci_respF_6$enq_1__SEL_6 =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_F_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_F_T_T_T ;
  assign MUX_wci_respF_6$enq_1__SEL_7 =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_F_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_T_F ;
  assign MUX_wci_respF_7$enq_1__SEL_6 =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_F_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_F_T_T_T ;
  assign MUX_wci_respF_7$enq_1__SEL_7 =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_T_F ;
  assign MUX_wci_respF_8$enq_1__SEL_6 =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_F_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_F_T_T_T ;
  assign MUX_wci_respF_8$enq_1__SEL_7 =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_T_F ;
  assign MUX_wci_respF_9$enq_1__SEL_6 =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_F_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T ;
  assign MUX_wci_respF_9$enq_1__SEL_7 =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_T_F ;
  assign MUX_wrkAct$write_1__SEL_1 =
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_F_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_F_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_F_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_F_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_F_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_F_F_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_F_F_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_F_F_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_T_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_T_F_F_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_T_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_T_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_T_F_F_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_T_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_T_T_T ;
  assign MUX_wrkAct$write_1__SEL_2 =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_F_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_F_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_F_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_F_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_F_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_F_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_F_F_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_F_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_F_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_F_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_F_F_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_F_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_F_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_F_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_F_F_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_F_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_F_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_F_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_T_F_F_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_T_F_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_T_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_T_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_T_F_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_T_F_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_T_T_T ;
  assign MUX_wrkAct$write_1__SEL_3 =
	     WILL_FIRE_RL_completeWorkerRead ||
	     WILL_FIRE_RL_completeWorkerWrite ;
  assign MUX_adminResp2F$enq_1__VAL_1 =
	     { cpReq[11:4] == 8'h30 || cpReq[11:4] == 8'h34 ||
	       cpReq[11:4] == 8'h38 ||
	       cpReq[11:4] == 8'h3C ||
	       cpReq[11:4] == 8'h40 ||
	       cpReq[11:4] == 8'h44 ||
	       cpReq[11:4] == 8'h48 ||
	       cpReq[11:4] == 8'h4C ||
	       cpReq[11:4] == 8'h50 ||
	       cpReq[11:4] == 8'h54 ||
	       cpReq[11:4] == 8'h7C ||
	       cpReq[11:4] == 8'h80 ||
	       cpReq[11:4] == 8'h84,
	       IF_cpReq_363_BITS_11_TO_4_366_EQ_0x30_595_THEN_ETC___d6177 } ;
  assign MUX_adminResp2F$enq_1__VAL_2 =
	     { 1'd1,
	       IF_cpReq_363_BITS_11_TO_4_366_EQ_0x30_595_THEN_ETC___d6177 } ;
  assign MUX_adminResp2F$enq_1__VAL_3 =
	     { cpReq[11:4] == 8'h50 || cpReq[11:4] == 8'h54 ||
	       cpReq[11:4] == 8'h7C ||
	       cpReq[11:4] == 8'h80 ||
	       cpReq[11:4] == 8'h84,
	       IF_cpReq_363_BITS_11_TO_4_366_EQ_0x30_595_THEN_ETC___d6177 } ;
  assign MUX_cpReq$write_1__VAL_4 =
	     cpReqF$D_OUT[58] ?
	       { (cpReqF$D_OUT[25:18] == 8'd0) ? 3'd2 : 3'd4,
		 24'hAAAAAA,
		 (cpReqF$D_OUT[25:18] == 8'd0) ?
		   2'd0 :
		   ((cpReqF$D_OUT[25:22] == 4'd0) ? 2'd1 : 2'd2),
		 cpReqF$D_OUT[33:26],
		 bAddr__h114303,
		 cpReqF$D_OUT[3:0] } :
	       { (cpReqF$D_OUT[57:50] == 8'd0) ?
		   5'd4 :
		   ((cpReqF$D_OUT[57:54] == 4'd0) ? 5'd13 : 5'd14),
		 cpReqF$D_OUT[31:0],
		 bAddr__h113843,
		 cpReqF$D_OUT[35:32] } ;
  assign MUX_cpRespF$enq_1__VAL_1 = { seqTag, crr_data__h76602 } ;
  assign MUX_cpRespF$enq_1__VAL_2 = { cpReq[35:28], rtnData__h113334 } ;
  assign MUX_readCntReg$write_1__VAL_2 = readCntReg + 32'd1 ;
  always@(wci_reqPend or wci_reqERR)
  begin
    case (wci_reqPend)
      2'd1: MUX_wci_reqERR$write_1__VAL_1 = { 1'd1, wci_reqERR[1:0] };
      2'd2:
	  MUX_wci_reqERR$write_1__VAL_1 =
	      { wci_reqERR[2], 1'd1, wci_reqERR[0] };
      default: MUX_wci_reqERR$write_1__VAL_1 = { wci_reqERR[2:1], 1'd1 };
    endcase
  end
  always@(wci_reqPend_1 or wci_reqERR_1)
  begin
    case (wci_reqPend_1)
      2'd1: MUX_wci_reqERR_1$write_1__VAL_1 = { 1'd1, wci_reqERR_1[1:0] };
      2'd2:
	  MUX_wci_reqERR_1$write_1__VAL_1 =
	      { wci_reqERR_1[2], 1'd1, wci_reqERR_1[0] };
      default: MUX_wci_reqERR_1$write_1__VAL_1 = { wci_reqERR_1[2:1], 1'd1 };
    endcase
  end
  always@(wci_reqPend_10 or wci_reqERR_10)
  begin
    case (wci_reqPend_10)
      2'd1: MUX_wci_reqERR_10$write_1__VAL_1 = { 1'd1, wci_reqERR_10[1:0] };
      2'd2:
	  MUX_wci_reqERR_10$write_1__VAL_1 =
	      { wci_reqERR_10[2], 1'd1, wci_reqERR_10[0] };
      default: MUX_wci_reqERR_10$write_1__VAL_1 =
		   { wci_reqERR_10[2:1], 1'd1 };
    endcase
  end
  always@(wci_reqPend_11 or wci_reqERR_11)
  begin
    case (wci_reqPend_11)
      2'd1: MUX_wci_reqERR_11$write_1__VAL_1 = { 1'd1, wci_reqERR_11[1:0] };
      2'd2:
	  MUX_wci_reqERR_11$write_1__VAL_1 =
	      { wci_reqERR_11[2], 1'd1, wci_reqERR_11[0] };
      default: MUX_wci_reqERR_11$write_1__VAL_1 =
		   { wci_reqERR_11[2:1], 1'd1 };
    endcase
  end
  always@(wci_reqPend_12 or wci_reqERR_12)
  begin
    case (wci_reqPend_12)
      2'd1: MUX_wci_reqERR_12$write_1__VAL_1 = { 1'd1, wci_reqERR_12[1:0] };
      2'd2:
	  MUX_wci_reqERR_12$write_1__VAL_1 =
	      { wci_reqERR_12[2], 1'd1, wci_reqERR_12[0] };
      default: MUX_wci_reqERR_12$write_1__VAL_1 =
		   { wci_reqERR_12[2:1], 1'd1 };
    endcase
  end
  always@(wci_reqPend_13 or wci_reqERR_13)
  begin
    case (wci_reqPend_13)
      2'd1: MUX_wci_reqERR_13$write_1__VAL_1 = { 1'd1, wci_reqERR_13[1:0] };
      2'd2:
	  MUX_wci_reqERR_13$write_1__VAL_1 =
	      { wci_reqERR_13[2], 1'd1, wci_reqERR_13[0] };
      default: MUX_wci_reqERR_13$write_1__VAL_1 =
		   { wci_reqERR_13[2:1], 1'd1 };
    endcase
  end
  always@(wci_reqPend_14 or wci_reqERR_14)
  begin
    case (wci_reqPend_14)
      2'd1: MUX_wci_reqERR_14$write_1__VAL_1 = { 1'd1, wci_reqERR_14[1:0] };
      2'd2:
	  MUX_wci_reqERR_14$write_1__VAL_1 =
	      { wci_reqERR_14[2], 1'd1, wci_reqERR_14[0] };
      default: MUX_wci_reqERR_14$write_1__VAL_1 =
		   { wci_reqERR_14[2:1], 1'd1 };
    endcase
  end
  always@(wci_reqPend_2 or wci_reqERR_2)
  begin
    case (wci_reqPend_2)
      2'd1: MUX_wci_reqERR_2$write_1__VAL_1 = { 1'd1, wci_reqERR_2[1:0] };
      2'd2:
	  MUX_wci_reqERR_2$write_1__VAL_1 =
	      { wci_reqERR_2[2], 1'd1, wci_reqERR_2[0] };
      default: MUX_wci_reqERR_2$write_1__VAL_1 = { wci_reqERR_2[2:1], 1'd1 };
    endcase
  end
  always@(wci_reqPend_3 or wci_reqERR_3)
  begin
    case (wci_reqPend_3)
      2'd1: MUX_wci_reqERR_3$write_1__VAL_1 = { 1'd1, wci_reqERR_3[1:0] };
      2'd2:
	  MUX_wci_reqERR_3$write_1__VAL_1 =
	      { wci_reqERR_3[2], 1'd1, wci_reqERR_3[0] };
      default: MUX_wci_reqERR_3$write_1__VAL_1 = { wci_reqERR_3[2:1], 1'd1 };
    endcase
  end
  always@(wci_reqPend_4 or wci_reqERR_4)
  begin
    case (wci_reqPend_4)
      2'd1: MUX_wci_reqERR_4$write_1__VAL_1 = { 1'd1, wci_reqERR_4[1:0] };
      2'd2:
	  MUX_wci_reqERR_4$write_1__VAL_1 =
	      { wci_reqERR_4[2], 1'd1, wci_reqERR_4[0] };
      default: MUX_wci_reqERR_4$write_1__VAL_1 = { wci_reqERR_4[2:1], 1'd1 };
    endcase
  end
  always@(wci_reqPend_5 or wci_reqERR_5)
  begin
    case (wci_reqPend_5)
      2'd1: MUX_wci_reqERR_5$write_1__VAL_1 = { 1'd1, wci_reqERR_5[1:0] };
      2'd2:
	  MUX_wci_reqERR_5$write_1__VAL_1 =
	      { wci_reqERR_5[2], 1'd1, wci_reqERR_5[0] };
      default: MUX_wci_reqERR_5$write_1__VAL_1 = { wci_reqERR_5[2:1], 1'd1 };
    endcase
  end
  always@(wci_reqPend_6 or wci_reqERR_6)
  begin
    case (wci_reqPend_6)
      2'd1: MUX_wci_reqERR_6$write_1__VAL_1 = { 1'd1, wci_reqERR_6[1:0] };
      2'd2:
	  MUX_wci_reqERR_6$write_1__VAL_1 =
	      { wci_reqERR_6[2], 1'd1, wci_reqERR_6[0] };
      default: MUX_wci_reqERR_6$write_1__VAL_1 = { wci_reqERR_6[2:1], 1'd1 };
    endcase
  end
  always@(wci_reqPend_7 or wci_reqERR_7)
  begin
    case (wci_reqPend_7)
      2'd1: MUX_wci_reqERR_7$write_1__VAL_1 = { 1'd1, wci_reqERR_7[1:0] };
      2'd2:
	  MUX_wci_reqERR_7$write_1__VAL_1 =
	      { wci_reqERR_7[2], 1'd1, wci_reqERR_7[0] };
      default: MUX_wci_reqERR_7$write_1__VAL_1 = { wci_reqERR_7[2:1], 1'd1 };
    endcase
  end
  always@(wci_reqPend_8 or wci_reqERR_8)
  begin
    case (wci_reqPend_8)
      2'd1: MUX_wci_reqERR_8$write_1__VAL_1 = { 1'd1, wci_reqERR_8[1:0] };
      2'd2:
	  MUX_wci_reqERR_8$write_1__VAL_1 =
	      { wci_reqERR_8[2], 1'd1, wci_reqERR_8[0] };
      default: MUX_wci_reqERR_8$write_1__VAL_1 = { wci_reqERR_8[2:1], 1'd1 };
    endcase
  end
  always@(wci_reqPend_9 or wci_reqERR_9)
  begin
    case (wci_reqPend_9)
      2'd1: MUX_wci_reqERR_9$write_1__VAL_1 = { 1'd1, wci_reqERR_9[1:0] };
      2'd2:
	  MUX_wci_reqERR_9$write_1__VAL_1 =
	      { wci_reqERR_9[2], 1'd1, wci_reqERR_9[0] };
      default: MUX_wci_reqERR_9$write_1__VAL_1 = { wci_reqERR_9[2:1], 1'd1 };
    endcase
  end
  always@(wci_reqPend or wci_reqFAIL)
  begin
    case (wci_reqPend)
      2'd1: MUX_wci_reqFAIL$write_1__VAL_1 = { 1'd1, wci_reqFAIL[1:0] };
      2'd2:
	  MUX_wci_reqFAIL$write_1__VAL_1 =
	      { wci_reqFAIL[2], 1'd1, wci_reqFAIL[0] };
      default: MUX_wci_reqFAIL$write_1__VAL_1 = { wci_reqFAIL[2:1], 1'd1 };
    endcase
  end
  always@(wci_reqPend_1 or wci_reqFAIL_1)
  begin
    case (wci_reqPend_1)
      2'd1: MUX_wci_reqFAIL_1$write_1__VAL_1 = { 1'd1, wci_reqFAIL_1[1:0] };
      2'd2:
	  MUX_wci_reqFAIL_1$write_1__VAL_1 =
	      { wci_reqFAIL_1[2], 1'd1, wci_reqFAIL_1[0] };
      default: MUX_wci_reqFAIL_1$write_1__VAL_1 =
		   { wci_reqFAIL_1[2:1], 1'd1 };
    endcase
  end
  always@(wci_reqPend_10 or wci_reqFAIL_10)
  begin
    case (wci_reqPend_10)
      2'd1: MUX_wci_reqFAIL_10$write_1__VAL_1 = { 1'd1, wci_reqFAIL_10[1:0] };
      2'd2:
	  MUX_wci_reqFAIL_10$write_1__VAL_1 =
	      { wci_reqFAIL_10[2], 1'd1, wci_reqFAIL_10[0] };
      default: MUX_wci_reqFAIL_10$write_1__VAL_1 =
		   { wci_reqFAIL_10[2:1], 1'd1 };
    endcase
  end
  always@(wci_reqPend_11 or wci_reqFAIL_11)
  begin
    case (wci_reqPend_11)
      2'd1: MUX_wci_reqFAIL_11$write_1__VAL_1 = { 1'd1, wci_reqFAIL_11[1:0] };
      2'd2:
	  MUX_wci_reqFAIL_11$write_1__VAL_1 =
	      { wci_reqFAIL_11[2], 1'd1, wci_reqFAIL_11[0] };
      default: MUX_wci_reqFAIL_11$write_1__VAL_1 =
		   { wci_reqFAIL_11[2:1], 1'd1 };
    endcase
  end
  always@(wci_reqPend_12 or wci_reqFAIL_12)
  begin
    case (wci_reqPend_12)
      2'd1: MUX_wci_reqFAIL_12$write_1__VAL_1 = { 1'd1, wci_reqFAIL_12[1:0] };
      2'd2:
	  MUX_wci_reqFAIL_12$write_1__VAL_1 =
	      { wci_reqFAIL_12[2], 1'd1, wci_reqFAIL_12[0] };
      default: MUX_wci_reqFAIL_12$write_1__VAL_1 =
		   { wci_reqFAIL_12[2:1], 1'd1 };
    endcase
  end
  always@(wci_reqPend_13 or wci_reqFAIL_13)
  begin
    case (wci_reqPend_13)
      2'd1: MUX_wci_reqFAIL_13$write_1__VAL_1 = { 1'd1, wci_reqFAIL_13[1:0] };
      2'd2:
	  MUX_wci_reqFAIL_13$write_1__VAL_1 =
	      { wci_reqFAIL_13[2], 1'd1, wci_reqFAIL_13[0] };
      default: MUX_wci_reqFAIL_13$write_1__VAL_1 =
		   { wci_reqFAIL_13[2:1], 1'd1 };
    endcase
  end
  always@(wci_reqPend_14 or wci_reqFAIL_14)
  begin
    case (wci_reqPend_14)
      2'd1: MUX_wci_reqFAIL_14$write_1__VAL_1 = { 1'd1, wci_reqFAIL_14[1:0] };
      2'd2:
	  MUX_wci_reqFAIL_14$write_1__VAL_1 =
	      { wci_reqFAIL_14[2], 1'd1, wci_reqFAIL_14[0] };
      default: MUX_wci_reqFAIL_14$write_1__VAL_1 =
		   { wci_reqFAIL_14[2:1], 1'd1 };
    endcase
  end
  always@(wci_reqPend_2 or wci_reqFAIL_2)
  begin
    case (wci_reqPend_2)
      2'd1: MUX_wci_reqFAIL_2$write_1__VAL_1 = { 1'd1, wci_reqFAIL_2[1:0] };
      2'd2:
	  MUX_wci_reqFAIL_2$write_1__VAL_1 =
	      { wci_reqFAIL_2[2], 1'd1, wci_reqFAIL_2[0] };
      default: MUX_wci_reqFAIL_2$write_1__VAL_1 =
		   { wci_reqFAIL_2[2:1], 1'd1 };
    endcase
  end
  always@(wci_reqPend_3 or wci_reqFAIL_3)
  begin
    case (wci_reqPend_3)
      2'd1: MUX_wci_reqFAIL_3$write_1__VAL_1 = { 1'd1, wci_reqFAIL_3[1:0] };
      2'd2:
	  MUX_wci_reqFAIL_3$write_1__VAL_1 =
	      { wci_reqFAIL_3[2], 1'd1, wci_reqFAIL_3[0] };
      default: MUX_wci_reqFAIL_3$write_1__VAL_1 =
		   { wci_reqFAIL_3[2:1], 1'd1 };
    endcase
  end
  always@(wci_reqPend_4 or wci_reqFAIL_4)
  begin
    case (wci_reqPend_4)
      2'd1: MUX_wci_reqFAIL_4$write_1__VAL_1 = { 1'd1, wci_reqFAIL_4[1:0] };
      2'd2:
	  MUX_wci_reqFAIL_4$write_1__VAL_1 =
	      { wci_reqFAIL_4[2], 1'd1, wci_reqFAIL_4[0] };
      default: MUX_wci_reqFAIL_4$write_1__VAL_1 =
		   { wci_reqFAIL_4[2:1], 1'd1 };
    endcase
  end
  always@(wci_reqPend_5 or wci_reqFAIL_5)
  begin
    case (wci_reqPend_5)
      2'd1: MUX_wci_reqFAIL_5$write_1__VAL_1 = { 1'd1, wci_reqFAIL_5[1:0] };
      2'd2:
	  MUX_wci_reqFAIL_5$write_1__VAL_1 =
	      { wci_reqFAIL_5[2], 1'd1, wci_reqFAIL_5[0] };
      default: MUX_wci_reqFAIL_5$write_1__VAL_1 =
		   { wci_reqFAIL_5[2:1], 1'd1 };
    endcase
  end
  always@(wci_reqPend_6 or wci_reqFAIL_6)
  begin
    case (wci_reqPend_6)
      2'd1: MUX_wci_reqFAIL_6$write_1__VAL_1 = { 1'd1, wci_reqFAIL_6[1:0] };
      2'd2:
	  MUX_wci_reqFAIL_6$write_1__VAL_1 =
	      { wci_reqFAIL_6[2], 1'd1, wci_reqFAIL_6[0] };
      default: MUX_wci_reqFAIL_6$write_1__VAL_1 =
		   { wci_reqFAIL_6[2:1], 1'd1 };
    endcase
  end
  always@(wci_reqPend_7 or wci_reqFAIL_7)
  begin
    case (wci_reqPend_7)
      2'd1: MUX_wci_reqFAIL_7$write_1__VAL_1 = { 1'd1, wci_reqFAIL_7[1:0] };
      2'd2:
	  MUX_wci_reqFAIL_7$write_1__VAL_1 =
	      { wci_reqFAIL_7[2], 1'd1, wci_reqFAIL_7[0] };
      default: MUX_wci_reqFAIL_7$write_1__VAL_1 =
		   { wci_reqFAIL_7[2:1], 1'd1 };
    endcase
  end
  always@(wci_reqPend_8 or wci_reqFAIL_8)
  begin
    case (wci_reqPend_8)
      2'd1: MUX_wci_reqFAIL_8$write_1__VAL_1 = { 1'd1, wci_reqFAIL_8[1:0] };
      2'd2:
	  MUX_wci_reqFAIL_8$write_1__VAL_1 =
	      { wci_reqFAIL_8[2], 1'd1, wci_reqFAIL_8[0] };
      default: MUX_wci_reqFAIL_8$write_1__VAL_1 =
		   { wci_reqFAIL_8[2:1], 1'd1 };
    endcase
  end
  always@(wci_reqPend_9 or wci_reqFAIL_9)
  begin
    case (wci_reqPend_9)
      2'd1: MUX_wci_reqFAIL_9$write_1__VAL_1 = { 1'd1, wci_reqFAIL_9[1:0] };
      2'd2:
	  MUX_wci_reqFAIL_9$write_1__VAL_1 =
	      { wci_reqFAIL_9[2], 1'd1, wci_reqFAIL_9[0] };
      default: MUX_wci_reqFAIL_9$write_1__VAL_1 =
		   { wci_reqFAIL_9[2:1], 1'd1 };
    endcase
  end
  assign MUX_wci_reqF_10_c_r$write_1__VAL_1 = wci_reqF_10_c_r + 1'd1 ;
  assign MUX_wci_reqF_10_c_r$write_1__VAL_2 = wci_reqF_10_c_r - 1'd1 ;
  always@(WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_T_T or
	  MUX_wci_reqF_10_x_wire$wset_1__VAL_1 or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T or
	  MUX_wci_reqF_10_x_wire$wset_1__VAL_2 or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T or
	  MUX_wci_reqF_10_x_wire$wset_1__VAL_3)
  begin
    case (1'b1) // synopsys parallel_case
      WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_T_T:
	  MUX_wci_reqF_10_q_0$write_1__VAL_1 =
	      MUX_wci_reqF_10_x_wire$wset_1__VAL_1;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T:
	  MUX_wci_reqF_10_q_0$write_1__VAL_1 =
	      MUX_wci_reqF_10_x_wire$wset_1__VAL_2;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T:
	  MUX_wci_reqF_10_q_0$write_1__VAL_1 =
	      MUX_wci_reqF_10_x_wire$wset_1__VAL_3;
      default: MUX_wci_reqF_10_q_0$write_1__VAL_1 =
		   72'hAAAAAAAAAAAAAAAAAA /* unspecified value */ ;
    endcase
  end
  assign MUX_wci_reqF_10_q_0$write_1__VAL_2 =
	     wci_reqF_10_c_r ?
	       MUX_wci_reqF_10_q_0$write_1__VAL_1 :
	       72'h0000000000AAAAAAAA ;
  assign MUX_wci_reqF_10_x_wire$wset_1__VAL_1 =
	     { 4'd3, cpReq[3:0], wciAddr__h78989, cpReq[59:28] } ;
  assign MUX_wci_reqF_10_x_wire$wset_1__VAL_2 =
	     { 4'd5, cpReq[3:0], wciAddr__h78989, 32'hAAAAAAAA } ;
  assign MUX_wci_reqF_10_x_wire$wset_1__VAL_3 =
	     { 8'd79, x_addr__h98551, 32'hAAAAAAAA } ;
  assign MUX_wci_reqF_11_c_r$write_1__VAL_1 = wci_reqF_11_c_r + 1'd1 ;
  assign MUX_wci_reqF_11_c_r$write_1__VAL_2 = wci_reqF_11_c_r - 1'd1 ;
  always@(WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_T_T or
	  MUX_wci_reqF_11_x_wire$wset_1__VAL_1 or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T or
	  MUX_wci_reqF_11_x_wire$wset_1__VAL_2 or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T or
	  MUX_wci_reqF_10_x_wire$wset_1__VAL_3)
  begin
    case (1'b1) // synopsys parallel_case
      WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_T_T:
	  MUX_wci_reqF_11_q_0$write_1__VAL_1 =
	      MUX_wci_reqF_11_x_wire$wset_1__VAL_1;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T:
	  MUX_wci_reqF_11_q_0$write_1__VAL_1 =
	      MUX_wci_reqF_11_x_wire$wset_1__VAL_2;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T:
	  MUX_wci_reqF_11_q_0$write_1__VAL_1 =
	      MUX_wci_reqF_10_x_wire$wset_1__VAL_3;
      default: MUX_wci_reqF_11_q_0$write_1__VAL_1 =
		   72'hAAAAAAAAAAAAAAAAAA /* unspecified value */ ;
    endcase
  end
  assign MUX_wci_reqF_11_q_0$write_1__VAL_2 =
	     wci_reqF_11_c_r ?
	       MUX_wci_reqF_11_q_0$write_1__VAL_1 :
	       72'h0000000000AAAAAAAA ;
  assign MUX_wci_reqF_11_x_wire$wset_1__VAL_1 =
	     { 4'd3, cpReq[3:0], wciAddr__h79055, cpReq[59:28] } ;
  assign MUX_wci_reqF_11_x_wire$wset_1__VAL_2 =
	     { 4'd5, cpReq[3:0], wciAddr__h79055, 32'hAAAAAAAA } ;
  assign MUX_wci_reqF_12_c_r$write_1__VAL_1 = wci_reqF_12_c_r + 1'd1 ;
  assign MUX_wci_reqF_12_c_r$write_1__VAL_2 = wci_reqF_12_c_r - 1'd1 ;
  always@(WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T or
	  MUX_wci_reqF_12_x_wire$wset_1__VAL_1 or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T or
	  MUX_wci_reqF_12_x_wire$wset_1__VAL_2 or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T or
	  MUX_wci_reqF_10_x_wire$wset_1__VAL_3)
  begin
    case (1'b1) // synopsys parallel_case
      WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T:
	  MUX_wci_reqF_12_q_0$write_1__VAL_1 =
	      MUX_wci_reqF_12_x_wire$wset_1__VAL_1;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T:
	  MUX_wci_reqF_12_q_0$write_1__VAL_1 =
	      MUX_wci_reqF_12_x_wire$wset_1__VAL_2;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T:
	  MUX_wci_reqF_12_q_0$write_1__VAL_1 =
	      MUX_wci_reqF_10_x_wire$wset_1__VAL_3;
      default: MUX_wci_reqF_12_q_0$write_1__VAL_1 =
		   72'hAAAAAAAAAAAAAAAAAA /* unspecified value */ ;
    endcase
  end
  assign MUX_wci_reqF_12_q_0$write_1__VAL_2 =
	     wci_reqF_12_c_r ?
	       MUX_wci_reqF_12_q_0$write_1__VAL_1 :
	       72'h0000000000AAAAAAAA ;
  assign MUX_wci_reqF_12_x_wire$wset_1__VAL_1 =
	     { 4'd3, cpReq[3:0], wciAddr__h79121, cpReq[59:28] } ;
  assign MUX_wci_reqF_12_x_wire$wset_1__VAL_2 =
	     { 4'd5, cpReq[3:0], wciAddr__h79121, 32'hAAAAAAAA } ;
  assign MUX_wci_reqF_13_c_r$write_1__VAL_1 = wci_reqF_13_c_r + 1'd1 ;
  assign MUX_wci_reqF_13_c_r$write_1__VAL_2 = wci_reqF_13_c_r - 1'd1 ;
  always@(WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T or
	  MUX_wci_reqF_13_x_wire$wset_1__VAL_1 or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T or
	  MUX_wci_reqF_13_x_wire$wset_1__VAL_2 or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T or
	  MUX_wci_reqF_10_x_wire$wset_1__VAL_3)
  begin
    case (1'b1) // synopsys parallel_case
      WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T:
	  MUX_wci_reqF_13_q_0$write_1__VAL_1 =
	      MUX_wci_reqF_13_x_wire$wset_1__VAL_1;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T:
	  MUX_wci_reqF_13_q_0$write_1__VAL_1 =
	      MUX_wci_reqF_13_x_wire$wset_1__VAL_2;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T:
	  MUX_wci_reqF_13_q_0$write_1__VAL_1 =
	      MUX_wci_reqF_10_x_wire$wset_1__VAL_3;
      default: MUX_wci_reqF_13_q_0$write_1__VAL_1 =
		   72'hAAAAAAAAAAAAAAAAAA /* unspecified value */ ;
    endcase
  end
  assign MUX_wci_reqF_13_q_0$write_1__VAL_2 =
	     wci_reqF_13_c_r ?
	       MUX_wci_reqF_13_q_0$write_1__VAL_1 :
	       72'h0000000000AAAAAAAA ;
  assign MUX_wci_reqF_13_x_wire$wset_1__VAL_1 =
	     { 4'd3, cpReq[3:0], wciAddr__h79187, cpReq[59:28] } ;
  assign MUX_wci_reqF_13_x_wire$wset_1__VAL_2 =
	     { 4'd5, cpReq[3:0], wciAddr__h79187, 32'hAAAAAAAA } ;
  assign MUX_wci_reqF_14_c_r$write_1__VAL_1 = wci_reqF_14_c_r + 1'd1 ;
  assign MUX_wci_reqF_14_c_r$write_1__VAL_2 = wci_reqF_14_c_r - 1'd1 ;
  always@(WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T or
	  MUX_wci_reqF_14_x_wire$wset_1__VAL_1 or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T or
	  MUX_wci_reqF_14_x_wire$wset_1__VAL_2 or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T or
	  MUX_wci_reqF_10_x_wire$wset_1__VAL_3)
  begin
    case (1'b1) // synopsys parallel_case
      WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T:
	  MUX_wci_reqF_14_q_0$write_1__VAL_1 =
	      MUX_wci_reqF_14_x_wire$wset_1__VAL_1;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T:
	  MUX_wci_reqF_14_q_0$write_1__VAL_1 =
	      MUX_wci_reqF_14_x_wire$wset_1__VAL_2;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T:
	  MUX_wci_reqF_14_q_0$write_1__VAL_1 =
	      MUX_wci_reqF_10_x_wire$wset_1__VAL_3;
      default: MUX_wci_reqF_14_q_0$write_1__VAL_1 =
		   72'hAAAAAAAAAAAAAAAAAA /* unspecified value */ ;
    endcase
  end
  assign MUX_wci_reqF_14_q_0$write_1__VAL_2 =
	     wci_reqF_14_c_r ?
	       MUX_wci_reqF_14_q_0$write_1__VAL_1 :
	       72'h0000000000AAAAAAAA ;
  assign MUX_wci_reqF_14_x_wire$wset_1__VAL_1 =
	     { 4'd3, cpReq[3:0], wciAddr__h79253, cpReq[59:28] } ;
  assign MUX_wci_reqF_14_x_wire$wset_1__VAL_2 =
	     { 4'd5, cpReq[3:0], wciAddr__h79253, 32'hAAAAAAAA } ;
  assign MUX_wci_reqF_1_c_r$write_1__VAL_1 = wci_reqF_1_c_r + 1'd1 ;
  assign MUX_wci_reqF_1_c_r$write_1__VAL_2 = wci_reqF_1_c_r - 1'd1 ;
  assign MUX_wci_reqF_1_q_0$write_1__VAL_1 =
	     wci_reqF_1_c_r ?
	       MUX_wci_reqF_1_q_0$write_1__VAL_2 :
	       72'h0000000000AAAAAAAA ;
  always@(WILL_FIRE_RL_cpDispatch_F_F_T_F_T_T_T or
	  MUX_wci_reqF_1_x_wire$wset_1__VAL_1 or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_T_T or
	  MUX_wci_reqF_1_x_wire$wset_1__VAL_2 or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_F_T_T or
	  MUX_wci_reqF_10_x_wire$wset_1__VAL_3)
  begin
    case (1'b1) // synopsys parallel_case
      WILL_FIRE_RL_cpDispatch_F_F_T_F_T_T_T:
	  MUX_wci_reqF_1_q_0$write_1__VAL_2 =
	      MUX_wci_reqF_1_x_wire$wset_1__VAL_1;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_T_T:
	  MUX_wci_reqF_1_q_0$write_1__VAL_2 =
	      MUX_wci_reqF_1_x_wire$wset_1__VAL_2;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_F_T_T:
	  MUX_wci_reqF_1_q_0$write_1__VAL_2 =
	      MUX_wci_reqF_10_x_wire$wset_1__VAL_3;
      default: MUX_wci_reqF_1_q_0$write_1__VAL_2 =
		   72'hAAAAAAAAAAAAAAAAAA /* unspecified value */ ;
    endcase
  end
  assign MUX_wci_reqF_1_x_wire$wset_1__VAL_1 =
	     { 4'd3, cpReq[3:0], wciAddr__h78395, cpReq[59:28] } ;
  assign MUX_wci_reqF_1_x_wire$wset_1__VAL_2 =
	     { 4'd5, cpReq[3:0], wciAddr__h78395, 32'hAAAAAAAA } ;
  assign MUX_wci_reqF_2_c_r$write_1__VAL_1 = wci_reqF_2_c_r + 1'd1 ;
  assign MUX_wci_reqF_2_c_r$write_1__VAL_2 = wci_reqF_2_c_r - 1'd1 ;
  assign MUX_wci_reqF_2_q_0$write_1__VAL_1 =
	     wci_reqF_2_c_r ?
	       MUX_wci_reqF_2_q_0$write_1__VAL_2 :
	       72'h0000000000AAAAAAAA ;
  always@(WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_T_T or
	  MUX_wci_reqF_2_x_wire$wset_1__VAL_1 or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_T_T or
	  MUX_wci_reqF_2_x_wire$wset_1__VAL_2 or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_F_T_T or
	  MUX_wci_reqF_10_x_wire$wset_1__VAL_3)
  begin
    case (1'b1) // synopsys parallel_case
      WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_T_T:
	  MUX_wci_reqF_2_q_0$write_1__VAL_2 =
	      MUX_wci_reqF_2_x_wire$wset_1__VAL_1;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_T_T:
	  MUX_wci_reqF_2_q_0$write_1__VAL_2 =
	      MUX_wci_reqF_2_x_wire$wset_1__VAL_2;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_F_T_T:
	  MUX_wci_reqF_2_q_0$write_1__VAL_2 =
	      MUX_wci_reqF_10_x_wire$wset_1__VAL_3;
      default: MUX_wci_reqF_2_q_0$write_1__VAL_2 =
		   72'hAAAAAAAAAAAAAAAAAA /* unspecified value */ ;
    endcase
  end
  assign MUX_wci_reqF_2_x_wire$wset_1__VAL_1 =
	     { 4'd3, cpReq[3:0], wciAddr__h78461, cpReq[59:28] } ;
  assign MUX_wci_reqF_2_x_wire$wset_1__VAL_2 =
	     { 4'd5, cpReq[3:0], wciAddr__h78461, 32'hAAAAAAAA } ;
  assign MUX_wci_reqF_3_c_r$write_1__VAL_1 = wci_reqF_3_c_r + 1'd1 ;
  assign MUX_wci_reqF_3_c_r$write_1__VAL_2 = wci_reqF_3_c_r - 1'd1 ;
  assign MUX_wci_reqF_3_q_0$write_1__VAL_1 =
	     wci_reqF_3_c_r ?
	       MUX_wci_reqF_3_q_0$write_1__VAL_2 :
	       72'h0000000000AAAAAAAA ;
  always@(WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_T_T or
	  MUX_wci_reqF_3_x_wire$wset_1__VAL_1 or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_T_T or
	  MUX_wci_reqF_3_x_wire$wset_1__VAL_2 or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_F_T_T or
	  MUX_wci_reqF_10_x_wire$wset_1__VAL_3)
  begin
    case (1'b1) // synopsys parallel_case
      WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_T_T:
	  MUX_wci_reqF_3_q_0$write_1__VAL_2 =
	      MUX_wci_reqF_3_x_wire$wset_1__VAL_1;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_T_T:
	  MUX_wci_reqF_3_q_0$write_1__VAL_2 =
	      MUX_wci_reqF_3_x_wire$wset_1__VAL_2;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_F_T_T:
	  MUX_wci_reqF_3_q_0$write_1__VAL_2 =
	      MUX_wci_reqF_10_x_wire$wset_1__VAL_3;
      default: MUX_wci_reqF_3_q_0$write_1__VAL_2 =
		   72'hAAAAAAAAAAAAAAAAAA /* unspecified value */ ;
    endcase
  end
  assign MUX_wci_reqF_3_x_wire$wset_1__VAL_1 =
	     { 4'd3, cpReq[3:0], wciAddr__h78527, cpReq[59:28] } ;
  assign MUX_wci_reqF_3_x_wire$wset_1__VAL_2 =
	     { 4'd5, cpReq[3:0], wciAddr__h78527, 32'hAAAAAAAA } ;
  assign MUX_wci_reqF_4_c_r$write_1__VAL_1 = wci_reqF_4_c_r + 1'd1 ;
  assign MUX_wci_reqF_4_c_r$write_1__VAL_2 = wci_reqF_4_c_r - 1'd1 ;
  assign MUX_wci_reqF_4_q_0$write_1__VAL_1 =
	     wci_reqF_4_c_r ?
	       MUX_wci_reqF_4_q_0$write_1__VAL_2 :
	       72'h0000000000AAAAAAAA ;
  always@(WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_T_T or
	  MUX_wci_reqF_4_x_wire$wset_1__VAL_1 or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_T_T or
	  MUX_wci_reqF_4_x_wire$wset_1__VAL_2 or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_F_T_T or
	  MUX_wci_reqF_10_x_wire$wset_1__VAL_3)
  begin
    case (1'b1) // synopsys parallel_case
      WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_T_T:
	  MUX_wci_reqF_4_q_0$write_1__VAL_2 =
	      MUX_wci_reqF_4_x_wire$wset_1__VAL_1;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_T_T:
	  MUX_wci_reqF_4_q_0$write_1__VAL_2 =
	      MUX_wci_reqF_4_x_wire$wset_1__VAL_2;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_F_T_T:
	  MUX_wci_reqF_4_q_0$write_1__VAL_2 =
	      MUX_wci_reqF_10_x_wire$wset_1__VAL_3;
      default: MUX_wci_reqF_4_q_0$write_1__VAL_2 =
		   72'hAAAAAAAAAAAAAAAAAA /* unspecified value */ ;
    endcase
  end
  assign MUX_wci_reqF_4_x_wire$wset_1__VAL_1 =
	     { 4'd3, cpReq[3:0], wciAddr__h78593, cpReq[59:28] } ;
  assign MUX_wci_reqF_4_x_wire$wset_1__VAL_2 =
	     { 4'd5, cpReq[3:0], wciAddr__h78593, 32'hAAAAAAAA } ;
  assign MUX_wci_reqF_5_c_r$write_1__VAL_1 = wci_reqF_5_c_r + 1'd1 ;
  assign MUX_wci_reqF_5_c_r$write_1__VAL_2 = wci_reqF_5_c_r - 1'd1 ;
  assign MUX_wci_reqF_5_q_0$write_1__VAL_1 =
	     wci_reqF_5_c_r ?
	       MUX_wci_reqF_5_q_0$write_1__VAL_2 :
	       72'h0000000000AAAAAAAA ;
  always@(WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_T_T or
	  MUX_wci_reqF_5_x_wire$wset_1__VAL_1 or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_T_T or
	  MUX_wci_reqF_5_x_wire$wset_1__VAL_2 or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_F_T_T or
	  MUX_wci_reqF_10_x_wire$wset_1__VAL_3)
  begin
    case (1'b1) // synopsys parallel_case
      WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_T_T:
	  MUX_wci_reqF_5_q_0$write_1__VAL_2 =
	      MUX_wci_reqF_5_x_wire$wset_1__VAL_1;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_T_T:
	  MUX_wci_reqF_5_q_0$write_1__VAL_2 =
	      MUX_wci_reqF_5_x_wire$wset_1__VAL_2;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_F_T_T:
	  MUX_wci_reqF_5_q_0$write_1__VAL_2 =
	      MUX_wci_reqF_10_x_wire$wset_1__VAL_3;
      default: MUX_wci_reqF_5_q_0$write_1__VAL_2 =
		   72'hAAAAAAAAAAAAAAAAAA /* unspecified value */ ;
    endcase
  end
  assign MUX_wci_reqF_5_x_wire$wset_1__VAL_1 =
	     { 4'd3, cpReq[3:0], wciAddr__h78659, cpReq[59:28] } ;
  assign MUX_wci_reqF_5_x_wire$wset_1__VAL_2 =
	     { 4'd5, cpReq[3:0], wciAddr__h78659, 32'hAAAAAAAA } ;
  assign MUX_wci_reqF_6_c_r$write_1__VAL_1 = wci_reqF_6_c_r + 1'd1 ;
  assign MUX_wci_reqF_6_c_r$write_1__VAL_2 = wci_reqF_6_c_r - 1'd1 ;
  assign MUX_wci_reqF_6_q_0$write_1__VAL_1 =
	     wci_reqF_6_c_r ?
	       MUX_wci_reqF_6_q_0$write_1__VAL_2 :
	       72'h0000000000AAAAAAAA ;
  always@(WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_T_T or
	  MUX_wci_reqF_6_x_wire$wset_1__VAL_1 or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_T_T or
	  MUX_wci_reqF_6_x_wire$wset_1__VAL_2 or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_F_T_T or
	  MUX_wci_reqF_10_x_wire$wset_1__VAL_3)
  begin
    case (1'b1) // synopsys parallel_case
      WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_T_T:
	  MUX_wci_reqF_6_q_0$write_1__VAL_2 =
	      MUX_wci_reqF_6_x_wire$wset_1__VAL_1;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_T_T:
	  MUX_wci_reqF_6_q_0$write_1__VAL_2 =
	      MUX_wci_reqF_6_x_wire$wset_1__VAL_2;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_F_T_T:
	  MUX_wci_reqF_6_q_0$write_1__VAL_2 =
	      MUX_wci_reqF_10_x_wire$wset_1__VAL_3;
      default: MUX_wci_reqF_6_q_0$write_1__VAL_2 =
		   72'hAAAAAAAAAAAAAAAAAA /* unspecified value */ ;
    endcase
  end
  assign MUX_wci_reqF_6_x_wire$wset_1__VAL_1 =
	     { 4'd3, cpReq[3:0], wciAddr__h78725, cpReq[59:28] } ;
  assign MUX_wci_reqF_6_x_wire$wset_1__VAL_2 =
	     { 4'd5, cpReq[3:0], wciAddr__h78725, 32'hAAAAAAAA } ;
  assign MUX_wci_reqF_7_c_r$write_1__VAL_1 = wci_reqF_7_c_r + 1'd1 ;
  assign MUX_wci_reqF_7_c_r$write_1__VAL_2 = wci_reqF_7_c_r - 1'd1 ;
  assign MUX_wci_reqF_7_q_0$write_1__VAL_1 =
	     wci_reqF_7_c_r ?
	       MUX_wci_reqF_7_q_0$write_1__VAL_2 :
	       72'h0000000000AAAAAAAA ;
  always@(WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_T_T or
	  MUX_wci_reqF_7_x_wire$wset_1__VAL_1 or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_T_T or
	  MUX_wci_reqF_7_x_wire$wset_1__VAL_2 or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T or
	  MUX_wci_reqF_10_x_wire$wset_1__VAL_3)
  begin
    case (1'b1) // synopsys parallel_case
      WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_T_T:
	  MUX_wci_reqF_7_q_0$write_1__VAL_2 =
	      MUX_wci_reqF_7_x_wire$wset_1__VAL_1;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_T_T:
	  MUX_wci_reqF_7_q_0$write_1__VAL_2 =
	      MUX_wci_reqF_7_x_wire$wset_1__VAL_2;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T:
	  MUX_wci_reqF_7_q_0$write_1__VAL_2 =
	      MUX_wci_reqF_10_x_wire$wset_1__VAL_3;
      default: MUX_wci_reqF_7_q_0$write_1__VAL_2 =
		   72'hAAAAAAAAAAAAAAAAAA /* unspecified value */ ;
    endcase
  end
  assign MUX_wci_reqF_7_x_wire$wset_1__VAL_1 =
	     { 4'd3, cpReq[3:0], wciAddr__h78791, cpReq[59:28] } ;
  assign MUX_wci_reqF_7_x_wire$wset_1__VAL_2 =
	     { 4'd5, cpReq[3:0], wciAddr__h78791, 32'hAAAAAAAA } ;
  assign MUX_wci_reqF_8_c_r$write_1__VAL_1 = wci_reqF_8_c_r + 1'd1 ;
  assign MUX_wci_reqF_8_c_r$write_1__VAL_2 = wci_reqF_8_c_r - 1'd1 ;
  assign MUX_wci_reqF_8_q_0$write_1__VAL_1 =
	     wci_reqF_8_c_r ?
	       MUX_wci_reqF_8_q_0$write_1__VAL_2 :
	       72'h0000000000AAAAAAAA ;
  always@(WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_T_T or
	  MUX_wci_reqF_8_x_wire$wset_1__VAL_1 or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T or
	  MUX_wci_reqF_8_x_wire$wset_1__VAL_2 or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T or
	  MUX_wci_reqF_10_x_wire$wset_1__VAL_3)
  begin
    case (1'b1) // synopsys parallel_case
      WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_T_T:
	  MUX_wci_reqF_8_q_0$write_1__VAL_2 =
	      MUX_wci_reqF_8_x_wire$wset_1__VAL_1;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T:
	  MUX_wci_reqF_8_q_0$write_1__VAL_2 =
	      MUX_wci_reqF_8_x_wire$wset_1__VAL_2;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T:
	  MUX_wci_reqF_8_q_0$write_1__VAL_2 =
	      MUX_wci_reqF_10_x_wire$wset_1__VAL_3;
      default: MUX_wci_reqF_8_q_0$write_1__VAL_2 =
		   72'hAAAAAAAAAAAAAAAAAA /* unspecified value */ ;
    endcase
  end
  assign MUX_wci_reqF_8_x_wire$wset_1__VAL_1 =
	     { 4'd3, cpReq[3:0], wciAddr__h78857, cpReq[59:28] } ;
  assign MUX_wci_reqF_8_x_wire$wset_1__VAL_2 =
	     { 4'd5, cpReq[3:0], wciAddr__h78857, 32'hAAAAAAAA } ;
  assign MUX_wci_reqF_9_c_r$write_1__VAL_1 = wci_reqF_9_c_r + 1'd1 ;
  assign MUX_wci_reqF_9_c_r$write_1__VAL_2 = wci_reqF_9_c_r - 1'd1 ;
  assign MUX_wci_reqF_9_q_0$write_1__VAL_1 =
	     wci_reqF_9_c_r ?
	       MUX_wci_reqF_9_q_0$write_1__VAL_2 :
	       72'h0000000000AAAAAAAA ;
  always@(WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_T_T or
	  MUX_wci_reqF_9_x_wire$wset_1__VAL_1 or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T or
	  MUX_wci_reqF_9_x_wire$wset_1__VAL_2 or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T or
	  MUX_wci_reqF_10_x_wire$wset_1__VAL_3)
  begin
    case (1'b1) // synopsys parallel_case
      WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_T_T:
	  MUX_wci_reqF_9_q_0$write_1__VAL_2 =
	      MUX_wci_reqF_9_x_wire$wset_1__VAL_1;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T:
	  MUX_wci_reqF_9_q_0$write_1__VAL_2 =
	      MUX_wci_reqF_9_x_wire$wset_1__VAL_2;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T:
	  MUX_wci_reqF_9_q_0$write_1__VAL_2 =
	      MUX_wci_reqF_10_x_wire$wset_1__VAL_3;
      default: MUX_wci_reqF_9_q_0$write_1__VAL_2 =
		   72'hAAAAAAAAAAAAAAAAAA /* unspecified value */ ;
    endcase
  end
  assign MUX_wci_reqF_9_x_wire$wset_1__VAL_1 =
	     { 4'd3, cpReq[3:0], wciAddr__h78923, cpReq[59:28] } ;
  assign MUX_wci_reqF_9_x_wire$wset_1__VAL_2 =
	     { 4'd5, cpReq[3:0], wciAddr__h78923, 32'hAAAAAAAA } ;
  assign MUX_wci_reqF_c_r$write_1__VAL_1 = wci_reqF_c_r + 1'd1 ;
  assign MUX_wci_reqF_c_r$write_1__VAL_2 = wci_reqF_c_r - 1'd1 ;
  assign MUX_wci_reqF_q_0$write_1__VAL_1 =
	     wci_reqF_c_r ?
	       MUX_wci_reqF_q_0$write_1__VAL_2 :
	       72'h0000000000AAAAAAAA ;
  always@(WILL_FIRE_RL_cpDispatch_F_F_T_T_T_T or
	  MUX_wci_reqF_x_wire$wset_1__VAL_1 or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_T_T_T or
	  MUX_wci_reqF_x_wire$wset_1__VAL_2 or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_T_F_T_T or
	  MUX_wci_reqF_10_x_wire$wset_1__VAL_3)
  begin
    case (1'b1) // synopsys parallel_case
      WILL_FIRE_RL_cpDispatch_F_F_T_T_T_T:
	  MUX_wci_reqF_q_0$write_1__VAL_2 = MUX_wci_reqF_x_wire$wset_1__VAL_1;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_T_T_T:
	  MUX_wci_reqF_q_0$write_1__VAL_2 = MUX_wci_reqF_x_wire$wset_1__VAL_2;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_T_F_T_T:
	  MUX_wci_reqF_q_0$write_1__VAL_2 =
	      MUX_wci_reqF_10_x_wire$wset_1__VAL_3;
      default: MUX_wci_reqF_q_0$write_1__VAL_2 =
		   72'hAAAAAAAAAAAAAAAAAA /* unspecified value */ ;
    endcase
  end
  assign MUX_wci_reqF_x_wire$wset_1__VAL_1 =
	     { 4'd3, cpReq[3:0], wciAddr__h78327, cpReq[59:28] } ;
  assign MUX_wci_reqF_x_wire$wset_1__VAL_2 =
	     { 4'd5, cpReq[3:0], wciAddr__h78327, 32'hAAAAAAAA } ;
  always@(wci_reqPend or wci_reqTO)
  begin
    case (wci_reqPend)
      2'd1: MUX_wci_reqTO$write_1__VAL_1 = { 1'd1, wci_reqTO[1:0] };
      2'd2:
	  MUX_wci_reqTO$write_1__VAL_1 = { wci_reqTO[2], 1'd1, wci_reqTO[0] };
      default: MUX_wci_reqTO$write_1__VAL_1 = { wci_reqTO[2:1], 1'd1 };
    endcase
  end
  always@(wci_reqPend_1 or wci_reqTO_1)
  begin
    case (wci_reqPend_1)
      2'd1: MUX_wci_reqTO_1$write_1__VAL_1 = { 1'd1, wci_reqTO_1[1:0] };
      2'd2:
	  MUX_wci_reqTO_1$write_1__VAL_1 =
	      { wci_reqTO_1[2], 1'd1, wci_reqTO_1[0] };
      default: MUX_wci_reqTO_1$write_1__VAL_1 = { wci_reqTO_1[2:1], 1'd1 };
    endcase
  end
  always@(wci_reqPend_10 or wci_reqTO_10)
  begin
    case (wci_reqPend_10)
      2'd1: MUX_wci_reqTO_10$write_1__VAL_1 = { 1'd1, wci_reqTO_10[1:0] };
      2'd2:
	  MUX_wci_reqTO_10$write_1__VAL_1 =
	      { wci_reqTO_10[2], 1'd1, wci_reqTO_10[0] };
      default: MUX_wci_reqTO_10$write_1__VAL_1 = { wci_reqTO_10[2:1], 1'd1 };
    endcase
  end
  always@(wci_reqPend_11 or wci_reqTO_11)
  begin
    case (wci_reqPend_11)
      2'd1: MUX_wci_reqTO_11$write_1__VAL_1 = { 1'd1, wci_reqTO_11[1:0] };
      2'd2:
	  MUX_wci_reqTO_11$write_1__VAL_1 =
	      { wci_reqTO_11[2], 1'd1, wci_reqTO_11[0] };
      default: MUX_wci_reqTO_11$write_1__VAL_1 = { wci_reqTO_11[2:1], 1'd1 };
    endcase
  end
  always@(wci_reqPend_12 or wci_reqTO_12)
  begin
    case (wci_reqPend_12)
      2'd1: MUX_wci_reqTO_12$write_1__VAL_1 = { 1'd1, wci_reqTO_12[1:0] };
      2'd2:
	  MUX_wci_reqTO_12$write_1__VAL_1 =
	      { wci_reqTO_12[2], 1'd1, wci_reqTO_12[0] };
      default: MUX_wci_reqTO_12$write_1__VAL_1 = { wci_reqTO_12[2:1], 1'd1 };
    endcase
  end
  always@(wci_reqPend_13 or wci_reqTO_13)
  begin
    case (wci_reqPend_13)
      2'd1: MUX_wci_reqTO_13$write_1__VAL_1 = { 1'd1, wci_reqTO_13[1:0] };
      2'd2:
	  MUX_wci_reqTO_13$write_1__VAL_1 =
	      { wci_reqTO_13[2], 1'd1, wci_reqTO_13[0] };
      default: MUX_wci_reqTO_13$write_1__VAL_1 = { wci_reqTO_13[2:1], 1'd1 };
    endcase
  end
  always@(wci_reqPend_14 or wci_reqTO_14)
  begin
    case (wci_reqPend_14)
      2'd1: MUX_wci_reqTO_14$write_1__VAL_1 = { 1'd1, wci_reqTO_14[1:0] };
      2'd2:
	  MUX_wci_reqTO_14$write_1__VAL_1 =
	      { wci_reqTO_14[2], 1'd1, wci_reqTO_14[0] };
      default: MUX_wci_reqTO_14$write_1__VAL_1 = { wci_reqTO_14[2:1], 1'd1 };
    endcase
  end
  always@(wci_reqPend_2 or wci_reqTO_2)
  begin
    case (wci_reqPend_2)
      2'd1: MUX_wci_reqTO_2$write_1__VAL_1 = { 1'd1, wci_reqTO_2[1:0] };
      2'd2:
	  MUX_wci_reqTO_2$write_1__VAL_1 =
	      { wci_reqTO_2[2], 1'd1, wci_reqTO_2[0] };
      default: MUX_wci_reqTO_2$write_1__VAL_1 = { wci_reqTO_2[2:1], 1'd1 };
    endcase
  end
  always@(wci_reqPend_3 or wci_reqTO_3)
  begin
    case (wci_reqPend_3)
      2'd1: MUX_wci_reqTO_3$write_1__VAL_1 = { 1'd1, wci_reqTO_3[1:0] };
      2'd2:
	  MUX_wci_reqTO_3$write_1__VAL_1 =
	      { wci_reqTO_3[2], 1'd1, wci_reqTO_3[0] };
      default: MUX_wci_reqTO_3$write_1__VAL_1 = { wci_reqTO_3[2:1], 1'd1 };
    endcase
  end
  always@(wci_reqPend_4 or wci_reqTO_4)
  begin
    case (wci_reqPend_4)
      2'd1: MUX_wci_reqTO_4$write_1__VAL_1 = { 1'd1, wci_reqTO_4[1:0] };
      2'd2:
	  MUX_wci_reqTO_4$write_1__VAL_1 =
	      { wci_reqTO_4[2], 1'd1, wci_reqTO_4[0] };
      default: MUX_wci_reqTO_4$write_1__VAL_1 = { wci_reqTO_4[2:1], 1'd1 };
    endcase
  end
  always@(wci_reqPend_5 or wci_reqTO_5)
  begin
    case (wci_reqPend_5)
      2'd1: MUX_wci_reqTO_5$write_1__VAL_1 = { 1'd1, wci_reqTO_5[1:0] };
      2'd2:
	  MUX_wci_reqTO_5$write_1__VAL_1 =
	      { wci_reqTO_5[2], 1'd1, wci_reqTO_5[0] };
      default: MUX_wci_reqTO_5$write_1__VAL_1 = { wci_reqTO_5[2:1], 1'd1 };
    endcase
  end
  always@(wci_reqPend_6 or wci_reqTO_6)
  begin
    case (wci_reqPend_6)
      2'd1: MUX_wci_reqTO_6$write_1__VAL_1 = { 1'd1, wci_reqTO_6[1:0] };
      2'd2:
	  MUX_wci_reqTO_6$write_1__VAL_1 =
	      { wci_reqTO_6[2], 1'd1, wci_reqTO_6[0] };
      default: MUX_wci_reqTO_6$write_1__VAL_1 = { wci_reqTO_6[2:1], 1'd1 };
    endcase
  end
  always@(wci_reqPend_7 or wci_reqTO_7)
  begin
    case (wci_reqPend_7)
      2'd1: MUX_wci_reqTO_7$write_1__VAL_1 = { 1'd1, wci_reqTO_7[1:0] };
      2'd2:
	  MUX_wci_reqTO_7$write_1__VAL_1 =
	      { wci_reqTO_7[2], 1'd1, wci_reqTO_7[0] };
      default: MUX_wci_reqTO_7$write_1__VAL_1 = { wci_reqTO_7[2:1], 1'd1 };
    endcase
  end
  always@(wci_reqPend_8 or wci_reqTO_8)
  begin
    case (wci_reqPend_8)
      2'd1: MUX_wci_reqTO_8$write_1__VAL_1 = { 1'd1, wci_reqTO_8[1:0] };
      2'd2:
	  MUX_wci_reqTO_8$write_1__VAL_1 =
	      { wci_reqTO_8[2], 1'd1, wci_reqTO_8[0] };
      default: MUX_wci_reqTO_8$write_1__VAL_1 = { wci_reqTO_8[2:1], 1'd1 };
    endcase
  end
  always@(wci_reqPend_9 or wci_reqTO_9)
  begin
    case (wci_reqPend_9)
      2'd1: MUX_wci_reqTO_9$write_1__VAL_1 = { 1'd1, wci_reqTO_9[1:0] };
      2'd2:
	  MUX_wci_reqTO_9$write_1__VAL_1 =
	      { wci_reqTO_9[2], 1'd1, wci_reqTO_9[0] };
      default: MUX_wci_reqTO_9$write_1__VAL_1 = { wci_reqTO_9[2:1], 1'd1 };
    endcase
  end
  assign MUX_wci_respF$enq_1__VAL_1 =
	     (wci_wciResponse$wget[33:32] == 2'd0) ?
	       34'h1C0DE4203 : // timeout
`ifdef not
	       wci_wciResponse$wget ;
`else
	      // If an OCP error response or OCP fail response, with something pending,
	      // Return the error code, whatever the op (config wrt, read, control op)
	      ((wci_wciResponse$wget[33:32] == 2'd3 || wci_wciResponse$wget[33:32] == 2'd2) &&
	       wci_reqPend != 2'd0 ? 34'h1C0DE4202 :
	       // This is success.  Return success code for ctlop or cfgwrt, but data for cfg read
	       (wci_reqPend == 2'd1 || wci_reqPend == 2'd3 ? 34'h1C0DE4201 : wci_wciResponse$wget));
`endif	       
  assign MUX_wci_respF$enq_1__VAL_2 = { 2'd1, wci_wStatus } ;
  assign MUX_wci_respF$enq_1__VAL_3 = { 2'd1, x_data__h104757 } ;
  assign MUX_wci_respF$enq_1__VAL_4 = { 2'd1, x_data__h104763 } ;
  assign MUX_wci_respF$enq_1__VAL_5 = { 22'd1048576, wci_pageWindow } ;
  assign MUX_wci_respF_1$enq_1__VAL_1 =
	     (wci_wciResponse_1$wget[33:32] == 2'd0) ?
	       34'h1C0DE4203 : 
`ifdef not
	       wci_wciResponse_1$wget ;
`else
	      // If an OCP error response or OCP fail response, with something pending,
	      // Return the error code, whatever the op (config wrt, read, control op)
	      ((wci_wciResponse_1$wget[33:32] == 2'd3 || wci_wciResponse_1$wget[33:32] == 2'd2) &&
	       wci_reqPend_1 != 2'd0 ? 34'h1C0DE4202 :
	       // This is success.  Return success code for ctlop or cfgwrt, but data for cfg read
	       (wci_reqPend_1 == 2'd1 || wci_reqPend_1 == 2'd3 ? 34'h1C0DE4201 : wci_wciResponse_1$wget));
`endif	       
  assign MUX_wci_respF_1$enq_1__VAL_2 = { 2'd1, wci_wStatus_1 } ;
  assign MUX_wci_respF_1$enq_1__VAL_3 = { 2'd1, x_data__h104810 } ;
  assign MUX_wci_respF_1$enq_1__VAL_4 = { 2'd1, x_data__h104816 } ;
  assign MUX_wci_respF_1$enq_1__VAL_5 = { 22'd1048576, wci_pageWindow_1 } ;
  assign MUX_wci_respF_10$enq_1__VAL_1 =
	     (wci_wciResponse_10$wget[33:32] == 2'd0) ?
	       34'h1C0DE4203 :
`ifdef not
	       wci_wciResponse_10$wget ;
`else
	      // If an OCP error response or OCP fail response, with something pending,
	      // Return the error code, whatever the op (config wrt, read, control op)
	      ((wci_wciResponse_10$wget[33:32] == 2'd3 || wci_wciResponse_10$wget[33:32] == 2'd2) &&
	       wci_reqPend_10 != 2'd0 ? 34'h1C0DE4202 :
	       // This is success.  Return success code for ctlop or cfgwrt, but data for cfg read
	       (wci_reqPend_10 == 2'd1 || wci_reqPend_10 == 2'd3 ? 34'h1C0DE4201 : wci_wciResponse_10$wget));
`endif	       
  assign MUX_wci_respF_10$enq_1__VAL_2 = { 2'd1, wci_wStatus_10 } ;
  assign MUX_wci_respF_10$enq_1__VAL_3 = { 2'd1, x_data__h105287 } ;
  assign MUX_wci_respF_10$enq_1__VAL_4 = { 2'd1, x_data__h105293 } ;
  assign MUX_wci_respF_10$enq_1__VAL_5 = { 22'd1048576, wci_pageWindow_10 } ;
  assign MUX_wci_respF_11$enq_1__VAL_1 =
	     (wci_wciResponse_11$wget[33:32] == 2'd0) ?
	       34'h1C0DE4203 :
`ifdef not
	       wci_wciResponse_11$wget ;
`else
	      // If an OCP error response or OCP fail response, with something pending,
	      // Return the error code, whatever the op (config wrt, read, control op)
	      ((wci_wciResponse_11$wget[33:32] == 2'd3 || wci_wciResponse_11$wget[33:32] == 2'd2) &&
	       wci_reqPend_11 != 2'd0 ? 34'h1C0DE4202 :
	       // This is success.  Return success code for ctlop or cfgwrt, but data for cfg read
	       (wci_reqPend_11 == 2'd1 || wci_reqPend_11 == 2'd3 ? 34'h1C0DE4201 : wci_wciResponse_11$wget));
`endif	       
  assign MUX_wci_respF_11$enq_1__VAL_2 = { 2'd1, wci_wStatus_11 } ;
  assign MUX_wci_respF_11$enq_1__VAL_3 = { 2'd1, x_data__h105340 } ;
  assign MUX_wci_respF_11$enq_1__VAL_4 = { 2'd1, x_data__h105346 } ;
  assign MUX_wci_respF_11$enq_1__VAL_5 = { 22'd1048576, wci_pageWindow_11 } ;
  assign MUX_wci_respF_12$enq_1__VAL_1 =
	     (wci_wciResponse_12$wget[33:32] == 2'd0) ?
	       34'h1C0DE4203 :
`ifdef not
	       wci_wciResponse_12$wget ;
`else
	      // If an OCP error response or OCP fail response, with something pending,
	      // Return the error code, whatever the op (config wrt, read, control op)
	      ((wci_wciResponse_12$wget[33:32] == 2'd3 || wci_wciResponse_12$wget[33:32] == 2'd2) &&
	       wci_reqPend_12 != 2'd0 ? 34'h1C0DE4202 :
	       // This is success.  Return success code for ctlop or cfgwrt, but data for cfg read
	       (wci_reqPend_12 == 2'd1 || wci_reqPend_12 == 2'd3 ? 34'h1C0DE4201 : wci_wciResponse_12$wget));
`endif	       
  assign MUX_wci_respF_12$enq_1__VAL_2 = { 2'd1, wci_wStatus_12 } ;
  assign MUX_wci_respF_12$enq_1__VAL_3 = { 2'd1, x_data__h105393 } ;
  assign MUX_wci_respF_12$enq_1__VAL_4 = { 2'd1, x_data__h105399 } ;
  assign MUX_wci_respF_12$enq_1__VAL_5 = { 22'd1048576, wci_pageWindow_12 } ;
  assign MUX_wci_respF_13$enq_1__VAL_1 =
	     (wci_wciResponse_13$wget[33:32] == 2'd0) ?
	       34'h1C0DE4203 :
`ifdef not
	       wci_wciResponse_13$wget ;
`else
	      // If an OCP error response or OCP fail response, with something pending,
	      // Return the error code, whatever the op (config wrt, read, control op)
	      ((wci_wciResponse_13$wget[33:32] == 2'd3 || wci_wciResponse_13$wget[33:32] == 2'd2) &&
	       wci_reqPend_13 != 2'd0 ? 34'h1C0DE4202 :
	       // This is success.  Return success code for ctlop or cfgwrt, but data for cfg read
	       (wci_reqPend_13 == 2'd1 || wci_reqPend_13 == 2'd3 ? 34'h1C0DE4201 : wci_wciResponse_13$wget));
`endif	       
  assign MUX_wci_respF_13$enq_1__VAL_2 = { 2'd1, wci_wStatus_13 } ;
  assign MUX_wci_respF_13$enq_1__VAL_3 = { 2'd1, x_data__h105446 } ;
  assign MUX_wci_respF_13$enq_1__VAL_4 = { 2'd1, x_data__h105452 } ;
  assign MUX_wci_respF_13$enq_1__VAL_5 = { 22'd1048576, wci_pageWindow_13 } ;
  assign MUX_wci_respF_14$enq_1__VAL_1 =
	     (wci_wciResponse_14$wget[33:32] == 2'd0) ?
	       34'h1C0DE4203 :
`ifdef not
	       wci_wciResponse_14$wget ;
`else
	      // If an OCP error response or OCP fail response, with something pending,
	      // Return the error code, whatever the op (config wrt, read, control op)
	      ((wci_wciResponse_14$wget[33:32] == 2'd3 || wci_wciResponse_14$wget[33:32] == 2'd2) &&
	       wci_reqPend_14 != 2'd0 ? 34'h1C0DE4202 :
	       // This is success.  Return success code for ctlop or cfgwrt, but data for cfg read
	       (wci_reqPend_14 == 2'd1 || wci_reqPend_14 == 2'd3 ? 34'h1C0DE4201 : wci_wciResponse_14$wget));
`endif	       
  assign MUX_wci_respF_14$enq_1__VAL_2 = { 2'd1, wci_wStatus_14 } ;
  assign MUX_wci_respF_14$enq_1__VAL_3 = { 2'd1, x_data__h105499 } ;
  assign MUX_wci_respF_14$enq_1__VAL_4 = { 2'd1, x_data__h105505 } ;
  assign MUX_wci_respF_14$enq_1__VAL_5 = { 22'd1048576, wci_pageWindow_14 } ;
  assign MUX_wci_respF_2$enq_1__VAL_1 =
	     (wci_wciResponse_2$wget[33:32] == 2'd0) ?
	       34'h1C0DE4203 :
`ifdef not
	       wci_wciResponse_2$wget ;
`else
	      // If an OCP error response or OCP fail response, with something pending,
	      // Return the error code, whatever the op (config wrt, read, control op)
	      ((wci_wciResponse_2$wget[33:32] == 2'd3 || wci_wciResponse_2$wget[33:32] == 2'd2) &&
	       wci_reqPend_2 != 2'd0 ? 34'h1C0DE4202 :
	       // This is success.  Return success code for ctlop or cfgwrt, but data for cfg read
	       (wci_reqPend_2 == 2'd1 || wci_reqPend_2 == 2'd3 ? 34'h1C0DE4201 : wci_wciResponse_2$wget));
`endif	       
  assign MUX_wci_respF_2$enq_1__VAL_2 = { 2'd1, wci_wStatus_2 } ;
  assign MUX_wci_respF_2$enq_1__VAL_3 = { 2'd1, x_data__h104863 } ;
  assign MUX_wci_respF_2$enq_1__VAL_4 = { 2'd1, x_data__h104869 } ;
  assign MUX_wci_respF_2$enq_1__VAL_5 = { 22'd1048576, wci_pageWindow_2 } ;
  assign MUX_wci_respF_3$enq_1__VAL_1 =
	     (wci_wciResponse_3$wget[33:32] == 2'd0) ?
	       34'h1C0DE4203 :
`ifdef not
	       wci_wciResponse_3$wget ;
`else
	      // If an OCP error response or OCP fail response, with something pending,
	      // Return the error code, whatever the op (config wrt, read, control op)
	      ((wci_wciResponse_3$wget[33:32] == 2'd3 || wci_wciResponse_3$wget[33:32] == 2'd2) &&
	       wci_reqPend_3 != 2'd0 ? 34'h1C0DE4202 :
	       // This is success.  Return success code for ctlop or cfgwrt, but data for cfg read
	       (wci_reqPend_3 == 2'd1 || wci_reqPend_3 == 2'd3 ? 34'h1C0DE4201 : wci_wciResponse_3$wget));
`endif	       
  assign MUX_wci_respF_3$enq_1__VAL_2 = { 2'd1, wci_wStatus_3 } ;
  assign MUX_wci_respF_3$enq_1__VAL_3 = { 2'd1, x_data__h104916 } ;
  assign MUX_wci_respF_3$enq_1__VAL_4 = { 2'd1, x_data__h104922 } ;
  assign MUX_wci_respF_3$enq_1__VAL_5 = { 22'd1048576, wci_pageWindow_3 } ;
  assign MUX_wci_respF_4$enq_1__VAL_1 =
	     (wci_wciResponse_4$wget[33:32] == 2'd0) ?
	       34'h1C0DE4203 :
`ifdef not
	       wci_wciResponse_4$wget ;
`else
	      // If an OCP error response or OCP fail response, with something pending,
	      // Return the error code, whatever the op (config wrt, read, control op)
	      ((wci_wciResponse_4$wget[33:32] == 2'd3 || wci_wciResponse_4$wget[33:32] == 2'd2) &&
	       wci_reqPend_4 != 2'd0 ? 34'h1C0DE4202 :
	       // This is success.  Return success code for ctlop or cfgwrt, but data for cfg read
	       (wci_reqPend_4 == 2'd1 || wci_reqPend_4 == 2'd3 ? 34'h1C0DE4201 : wci_wciResponse_4$wget));
`endif	       
  assign MUX_wci_respF_4$enq_1__VAL_2 = { 2'd1, wci_wStatus_4 } ;
  assign MUX_wci_respF_4$enq_1__VAL_3 = { 2'd1, x_data__h104969 } ;
  assign MUX_wci_respF_4$enq_1__VAL_4 = { 2'd1, x_data__h104975 } ;
  assign MUX_wci_respF_4$enq_1__VAL_5 = { 22'd1048576, wci_pageWindow_4 } ;
  assign MUX_wci_respF_5$enq_1__VAL_1 =
	     (wci_wciResponse_5$wget[33:32] == 2'd0) ?
	       34'h1C0DE4203 :
`ifdef not
	       wci_wciResponse_5$wget ;
`else
	      // If an OCP error response or OCP fail response, with something pending,
	      // Return the error code, whatever the op (config wrt, read, control op)
	      ((wci_wciResponse_5$wget[33:32] == 2'd3 || wci_wciResponse_5$wget[33:32] == 2'd2) &&
	       wci_reqPend_5 != 2'd0 ? 34'h1C0DE4202 :
	       // This is success.  Return success code for ctlop or cfgwrt, but data for cfg read
	       (wci_reqPend_5 == 2'd1 || wci_reqPend_5 == 2'd3 ? 34'h1C0DE4201 : wci_wciResponse_5$wget));
`endif	       
  assign MUX_wci_respF_5$enq_1__VAL_2 = { 2'd1, wci_wStatus_5 } ;
  assign MUX_wci_respF_5$enq_1__VAL_3 = { 2'd1, x_data__h105022 } ;
  assign MUX_wci_respF_5$enq_1__VAL_4 = { 2'd1, x_data__h105028 } ;
  assign MUX_wci_respF_5$enq_1__VAL_5 = { 22'd1048576, wci_pageWindow_5 } ;
  assign MUX_wci_respF_6$enq_1__VAL_1 =
	     (wci_wciResponse_6$wget[33:32] == 2'd0) ?
	       34'h1C0DE4203 :
`ifdef not
	       wci_wciResponse_6$wget ;
`else
	      // If an OCP error response or OCP fail response, with something pending,
	      // Return the error code, whatever the op (config wrt, read, control op)
	      ((wci_wciResponse_6$wget[33:32] == 2'd3 || wci_wciResponse_6$wget[33:32] == 2'd2) &&
	       wci_reqPend_6 != 2'd0 ? 34'h1C0DE4202 :
	       // This is success.  Return success code for ctlop or cfgwrt, but data for cfg read
	       (wci_reqPend_6 == 2'd1 || wci_reqPend_6 == 2'd3 ? 34'h1C0DE4201 : wci_wciResponse_6$wget));
`endif	       
  assign MUX_wci_respF_6$enq_1__VAL_2 = { 2'd1, wci_wStatus_6 } ;
  assign MUX_wci_respF_6$enq_1__VAL_3 = { 2'd1, x_data__h105075 } ;
  assign MUX_wci_respF_6$enq_1__VAL_4 = { 2'd1, x_data__h105081 } ;
  assign MUX_wci_respF_6$enq_1__VAL_5 = { 22'd1048576, wci_pageWindow_6 } ;
  assign MUX_wci_respF_7$enq_1__VAL_1 =
	     (wci_wciResponse_7$wget[33:32] == 2'd0) ?
	       34'h1C0DE4203 :
`ifdef not
	       wci_wciResponse_7$wget ;
`else
	      // If an OCP error response or OCP fail response, with something pending,
	      // Return the error code, whatever the op (config wrt, read, control op)
	      ((wci_wciResponse_7$wget[33:32] == 2'd3 || wci_wciResponse_7$wget[33:32] == 2'd2) &&
	       wci_reqPend_7 != 2'd0 ? 34'h1C0DE4202 :
	       // This is success.  Return success code for ctlop or cfgwrt, but data for cfg read
	       (wci_reqPend_7 == 2'd1 || wci_reqPend_7 == 2'd3 ? 34'h1C0DE4201 : wci_wciResponse_7$wget));
`endif	       
  assign MUX_wci_respF_7$enq_1__VAL_2 = { 2'd1, wci_wStatus_7 } ;
  assign MUX_wci_respF_7$enq_1__VAL_3 = { 2'd1, x_data__h105128 } ;
  assign MUX_wci_respF_7$enq_1__VAL_4 = { 2'd1, x_data__h105134 } ;
  assign MUX_wci_respF_7$enq_1__VAL_5 = { 22'd1048576, wci_pageWindow_7 } ;
  assign MUX_wci_respF_8$enq_1__VAL_1 =
	     (wci_wciResponse_8$wget[33:32] == 2'd0) ?
	       34'h1C0DE4203 :
`ifdef not
	       wci_wciResponse_8$wget ;
`else
	      // If an OCP error response or OCP fail response, with something pending,
	      // Return the error code, whatever the op (config wrt, read, control op)
	      ((wci_wciResponse_8$wget[33:32] == 2'd3 || wci_wciResponse_8$wget[33:32] == 2'd2) &&
	       wci_reqPend_8 != 2'd0 ? 34'h1C0DE4202 :
	       // This is success.  Return success code for ctlop or cfgwrt, but data for cfg read
	       (wci_reqPend_8 == 2'd1 || wci_reqPend_8 == 2'd3 ? 34'h1C0DE4201 : wci_wciResponse_8$wget));
`endif	       
  assign MUX_wci_respF_8$enq_1__VAL_2 = { 2'd1, wci_wStatus_8 } ;
  assign MUX_wci_respF_8$enq_1__VAL_3 = { 2'd1, x_data__h105181 } ;
  assign MUX_wci_respF_8$enq_1__VAL_4 = { 2'd1, x_data__h105187 } ;
  assign MUX_wci_respF_8$enq_1__VAL_5 = { 22'd1048576, wci_pageWindow_8 } ;
  assign MUX_wci_respF_9$enq_1__VAL_1 =
	     (wci_wciResponse_9$wget[33:32] == 2'd0) ?
	       34'h1C0DE4203 :
`ifdef not
	       wci_wciResponse_9$wget ;
`else
	      // If an OCP error response or OCP fail response, with something pending,
	      // Return the error code, whatever the op (config wrt, read, control op)
	      ((wci_wciResponse_9$wget[33:32] == 2'd3 || wci_wciResponse_9$wget[33:32] == 2'd2) &&
	       wci_reqPend_9 != 2'd0 ? 34'h1C0DE4202 :
	       // This is success.  Return success code for ctlop or cfgwrt, but data for cfg read
	       (wci_reqPend_9 == 2'd1 || wci_reqPend_9 == 2'd3 ? 34'h1C0DE4201 : wci_wciResponse_9$wget));
`endif	       
  assign MUX_wci_respF_9$enq_1__VAL_2 = { 2'd1, wci_wStatus_9 } ;
  assign MUX_wci_respF_9$enq_1__VAL_3 = { 2'd1, x_data__h105234 } ;
  assign MUX_wci_respF_9$enq_1__VAL_4 = { 2'd1, x_data__h105240 } ;
  assign MUX_wci_respF_9$enq_1__VAL_5 = { 22'd1048576, wci_pageWindow_9 } ;
  assign MUX_wci_respTimr$write_1__VAL_2 =
	     (wci_wciResponse$wget[33:32] == 2'd0) ?
	       (wci_respTimr_28_ULT_1_SL_wci_wTimeout_29_30___d5879 ?
		  x__h11924 :
		  32'd0) :
	       32'd0 ;
  assign MUX_wci_respTimr_1$write_1__VAL_2 =
	     (wci_wciResponse_1$wget[33:32] == 2'd0) ?
	       (wci_respTimr_1_68_ULT_1_SL_wci_wTimeout_1_69_70___d5880 ?
		  x__h16367 :
		  32'd0) :
	       32'd0 ;
  assign MUX_wci_respTimr_10$write_1__VAL_2 =
	     (wci_wciResponse_10$wget[33:32] == 2'd0) ?
	       (wci_respTimr_10_628_ULT_1_SL_wci_wTimeout_10_6_ETC___d5889 ?
		  x__h56327 :
		  32'd0) :
	       32'd0 ;
  assign MUX_wci_respTimr_11$write_1__VAL_2 =
	     (wci_wciResponse_11$wget[33:32] == 2'd0) ?
	       (wci_respTimr_11_768_ULT_1_SL_wci_wTimeout_11_7_ETC___d5890 ?
		  x__h60767 :
		  32'd0) :
	       32'd0 ;
  assign MUX_wci_respTimr_12$write_1__VAL_2 =
	     (wci_wciResponse_12$wget[33:32] == 2'd0) ?
	       (wci_respTimr_12_908_ULT_1_SL_wci_wTimeout_12_9_ETC___d5891 ?
		  x__h65207 :
		  32'd0) :
	       32'd0 ;
  assign MUX_wci_respTimr_13$write_1__VAL_2 =
	     (wci_wciResponse_13$wget[33:32] == 2'd0) ?
	       (wci_respTimr_13_048_ULT_1_SL_wci_wTimeout_13_0_ETC___d5892 ?
		  x__h69647 :
		  32'd0) :
	       32'd0 ;
  assign MUX_wci_respTimr_14$write_1__VAL_2 =
	     (wci_wciResponse_14$wget[33:32] == 2'd0) ?
	       (wci_respTimr_14_188_ULT_1_SL_wci_wTimeout_14_1_ETC___d5893 ?
		  x__h74087 :
		  32'd0) :
	       32'd0 ;
  assign MUX_wci_respTimr_2$write_1__VAL_2 =
	     (wci_wciResponse_2$wget[33:32] == 2'd0) ?
	       (wci_respTimr_2_08_ULT_1_SL_wci_wTimeout_2_09_10___d5881 ?
		  x__h20807 :
		  32'd0) :
	       32'd0 ;
  assign MUX_wci_respTimr_3$write_1__VAL_2 =
	     (wci_wciResponse_3$wget[33:32] == 2'd0) ?
	       (wci_respTimr_3_48_ULT_1_SL_wci_wTimeout_3_49_50___d5882 ?
		  x__h25247 :
		  32'd0) :
	       32'd0 ;
  assign MUX_wci_respTimr_4$write_1__VAL_2 =
	     (wci_wciResponse_4$wget[33:32] == 2'd0) ?
	       (wci_respTimr_4_88_ULT_1_SL_wci_wTimeout_4_89_90___d5883 ?
		  x__h29687 :
		  32'd0) :
	       32'd0 ;
  assign MUX_wci_respTimr_5$write_1__VAL_2 =
	     (wci_wciResponse_5$wget[33:32] == 2'd0) ?
	       (wci_respTimr_5_28_ULT_1_SL_wci_wTimeout_5_29_30___d5884 ?
		  x__h34127 :
		  32'd0) :
	       32'd0 ;
  assign MUX_wci_respTimr_6$write_1__VAL_2 =
	     (wci_wciResponse_6$wget[33:32] == 2'd0) ?
	       (wci_respTimr_6_068_ULT_1_SL_wci_wTimeout_6_069_ETC___d5885 ?
		  x__h38567 :
		  32'd0) :
	       32'd0 ;
  assign MUX_wci_respTimr_7$write_1__VAL_2 =
	     (wci_wciResponse_7$wget[33:32] == 2'd0) ?
	       (wci_respTimr_7_208_ULT_1_SL_wci_wTimeout_7_209_ETC___d5886 ?
		  x__h43007 :
		  32'd0) :
	       32'd0 ;
  assign MUX_wci_respTimr_8$write_1__VAL_2 =
	     (wci_wciResponse_8$wget[33:32] == 2'd0) ?
	       (wci_respTimr_8_348_ULT_1_SL_wci_wTimeout_8_349_ETC___d5887 ?
		  x__h47447 :
		  32'd0) :
	       32'd0 ;
  assign MUX_wci_respTimr_9$write_1__VAL_2 =
	     (wci_wciResponse_9$wget[33:32] == 2'd0) ?
	       (wci_respTimr_9_488_ULT_1_SL_wci_wTimeout_9_489_ETC___d5888 ?
		  x__h51887 :
		  32'd0) :
	       32'd0 ;

  // inlined wires
  assign warmResetP_1$wget = cpReq[59:28] == 32'hC0DEFFFF ;
  assign warmResetP_1$whas = WILL_FIRE_RL_cpDispatch_T_F_F_F_T ;
`ifdef not
  assign timeServ_jamFrac_1$wget = 1'd1 ;
  assign timeServ_jamFrac_1$whas =
	     timeServ_setRefF$dEMPTY_N && !timeServ_ppsOK ;
  assign timeServ_jamFracVal_1$wget = x__h3700 ;
  assign timeServ_jamFracVal_1$whas = timeServ_jamFrac_1$whas ;
  assign deviceDNA$wget = { 7'd0, dna_sr } ;
  assign deviceDNA$whas = dna_cnt == 7'd127 ;
  assign devDNAV$wget =
	     (dna_cnt == 7'd127) ? deviceDNA$wget : 64'h0BADC0DE0BADC0DE ;
  assign devDNAV$whas = 1'd1 ;
  assign rom_serverAdapter_outData_enqData$wget = rom_memory$DO ;
  assign rom_serverAdapter_outData_enqData$whas =
	     (!rom_serverAdapter_s1[0] ||
	      rom_serverAdapter_outDataCore$FULL_N) &&
	     rom_serverAdapter_s1[1] &&
	     rom_serverAdapter_s1[0] ;
  assign rom_serverAdapter_outData_outData$wget =
	     rom_serverAdapter_outDataCore$EMPTY_N ?
	       rom_serverAdapter_outDataCore$D_OUT :
	       rom_memory$DO ;
  assign rom_serverAdapter_outData_outData$whas =
	     rom_serverAdapter_outDataCore$EMPTY_N ||
	     !rom_serverAdapter_outDataCore$EMPTY_N &&
	     rom_serverAdapter_outData_enqData$whas ;
  assign rom_serverAdapter_cnt_1$wget = 3'd1 ;
  assign rom_serverAdapter_cnt_1$whas =
	     WILL_FIRE_RL_rom_serverAdapter_stageReadResponseAlways ;
  assign rom_serverAdapter_cnt_2$wget = 3'd7 ;
  assign rom_serverAdapter_cnt_2$whas =
	     rom_serverAdapter_outData_deqCalled$whas ;
  assign rom_serverAdapter_cnt_3$wget = 3'h0 ;
  assign rom_serverAdapter_cnt_3$whas = 1'b0 ;
  assign rom_serverAdapter_writeWithResp$wget = 2'd0 ;
  assign rom_serverAdapter_writeWithResp$whas =
	     WILL_FIRE_RL_rom_serverAdapter_stageReadResponseAlways ;
  assign rom_serverAdapter_s1_1$wget = 2'd3 ;
  assign rom_serverAdapter_s1_1$whas =
	     WILL_FIRE_RL_rom_serverAdapter_stageReadResponseAlways ;
  assign dna_rdReg_1$wget = 1'd1 ;
  assign dna_rdReg_1$whas = dna_cnt == 7'd1 || dna_cnt == 7'd2 ;
  assign dna_shftReg_1$wget = 1'd1 ;
  assign dna_shftReg_1$whas = dna_cnt >= 7'd3 && dna_cnt <= 7'd116 ;
  assign uuidV$wget = uuid_arg ;
  assign uuidV$whas = 1'd1 ;
  assign rom_memory$DO = rom_data;
  assign rom_addr = rom_memory$ADDR;
  assign rom_en = rom_memory$EN;
`endif
  assign wci_reqF_x_wire$wget = MUX_wci_reqF_q_0$write_1__VAL_2 ;
  assign wci_reqF_x_wire$whas =
	     WILL_FIRE_RL_cpDispatch_F_F_T_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_T_F_T_T ;
  assign wci_wciResponse$wget = { wci_Vm_0_SResp, wci_Vm_0_SData } ;
  assign wci_wciResponse$whas = 1'd1 ;
  assign wci_sfCapSet_1$wget = wci_Vm_0_SFlag[0] ;
  assign wci_sfCapSet_1$whas = 1'd1 ;
  assign wci_sfCapClear_1$wget = 1'd1 ;
  assign wci_sfCapClear_1$whas =
	     WILL_FIRE_RL_cpDispatch_F_F_T_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_T_F_F_T_T_T ;
  assign wci_reqF_1_x_wire$wget = MUX_wci_reqF_1_q_0$write_1__VAL_2 ;
  assign wci_reqF_1_x_wire$whas =
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_F_T_T ;
  assign wci_wciResponse_1$wget = { wci_Vm_1_SResp, wci_Vm_1_SData } ;
  assign wci_wciResponse_1$whas = 1'd1 ;
  assign wci_sfCapSet_1_2$wget = wci_Vm_1_SFlag[0] ;
  assign wci_sfCapSet_1_2$whas = 1'd1 ;
  assign wci_sfCapClear_1_2$wget = 1'd1 ;
  assign wci_sfCapClear_1_2$whas =
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_T_F_F_T_T_T ;
  assign wci_reqF_2_x_wire$wget = MUX_wci_reqF_2_q_0$write_1__VAL_2 ;
  assign wci_reqF_2_x_wire$whas =
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_F_T_T ;
  assign wci_wciResponse_2$wget = { wci_Vm_2_SResp, wci_Vm_2_SData } ;
  assign wci_wciResponse_2$whas = 1'd1 ;
  assign wci_sfCapSet_2_1$wget = wci_Vm_2_SFlag[0] ;
  assign wci_sfCapSet_2_1$whas = 1'd1 ;
  assign wci_sfCapClear_2_1$wget = 1'd1 ;
  assign wci_sfCapClear_2_1$whas =
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_F_F_T_T_T ;
  assign wci_reqF_3_x_wire$wget = MUX_wci_reqF_3_q_0$write_1__VAL_2 ;
  assign wci_reqF_3_x_wire$whas =
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_F_T_T ;
  assign wci_wciResponse_3$wget = { wci_Vm_3_SResp, wci_Vm_3_SData } ;
  assign wci_wciResponse_3$whas = 1'd1 ;
  assign wci_sfCapSet_3_1$wget = wci_Vm_3_SFlag[0] ;
  assign wci_sfCapSet_3_1$whas = 1'd1 ;
  assign wci_sfCapClear_3_1$wget = 1'd1 ;
  assign wci_sfCapClear_3_1$whas =
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_F_F_T_T_T ;
  assign wci_reqF_4_x_wire$wget = MUX_wci_reqF_4_q_0$write_1__VAL_2 ;
  assign wci_reqF_4_x_wire$whas =
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_F_T_T ;
  assign wci_wciResponse_4$wget = { wci_Vm_4_SResp, wci_Vm_4_SData } ;
  assign wci_wciResponse_4$whas = 1'd1 ;
  assign wci_sfCapSet_4_1$wget = wci_Vm_4_SFlag[0] ;
  assign wci_sfCapSet_4_1$whas = 1'd1 ;
  assign wci_sfCapClear_4_1$wget = 1'd1 ;
  assign wci_sfCapClear_4_1$whas =
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_F_F_T_T_T ;
  assign wci_reqF_5_x_wire$wget = MUX_wci_reqF_5_q_0$write_1__VAL_2 ;
  assign wci_reqF_5_x_wire$whas =
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_F_T_T ;
  assign wci_wciResponse_5$wget = { wci_Vm_5_SResp, wci_Vm_5_SData } ;
  assign wci_wciResponse_5$whas = 1'd1 ;
  assign wci_sfCapSet_5_1$wget = wci_Vm_5_SFlag[0] ;
  assign wci_sfCapSet_5_1$whas = 1'd1 ;
  assign wci_sfCapClear_5_1$wget = 1'd1 ;
  assign wci_sfCapClear_5_1$whas =
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_F_T_T_T ;
  assign wci_reqF_6_x_wire$wget = MUX_wci_reqF_6_q_0$write_1__VAL_2 ;
  assign wci_reqF_6_x_wire$whas =
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_F_T_T ;
  assign wci_wciResponse_6$wget = { wci_Vm_6_SResp, wci_Vm_6_SData } ;
  assign wci_wciResponse_6$whas = 1'd1 ;
  assign wci_sfCapSet_6_1$wget = wci_Vm_6_SFlag[0] ;
  assign wci_sfCapSet_6_1$whas = 1'd1 ;
  assign wci_sfCapClear_6_1$wget = 1'd1 ;
  assign wci_sfCapClear_6_1$whas =
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_F_T_T_T ;
  assign wci_reqF_7_x_wire$wget = MUX_wci_reqF_7_q_0$write_1__VAL_2 ;
  assign wci_reqF_7_x_wire$whas =
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T ;
  assign wci_wciResponse_7$wget = { wci_Vm_7_SResp, wci_Vm_7_SData } ;
  assign wci_wciResponse_7$whas = 1'd1 ;
  assign wci_sfCapSet_7_1$wget = wci_Vm_7_SFlag[0] ;
  assign wci_sfCapSet_7_1$whas = 1'd1 ;
  assign wci_sfCapClear_7_1$wget = 1'd1 ;
  assign wci_sfCapClear_7_1$whas =
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_F_T_T_T ;
  assign wci_reqF_8_x_wire$wget = MUX_wci_reqF_8_q_0$write_1__VAL_2 ;
  assign wci_reqF_8_x_wire$whas =
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T ;
  assign wci_wciResponse_8$wget = { wci_Vm_8_SResp, wci_Vm_8_SData } ;
  assign wci_wciResponse_8$whas = 1'd1 ;
  assign wci_sfCapSet_8_1$wget = wci_Vm_8_SFlag[0] ;
  assign wci_sfCapSet_8_1$whas = 1'd1 ;
  assign wci_sfCapClear_8_1$wget = 1'd1 ;
  assign wci_sfCapClear_8_1$whas =
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_F_T_T_T ;
  assign wci_reqF_9_x_wire$wget = MUX_wci_reqF_9_q_0$write_1__VAL_2 ;
  assign wci_reqF_9_x_wire$whas =
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T ;
  assign wci_wciResponse_9$wget = { wci_Vm_9_SResp, wci_Vm_9_SData } ;
  assign wci_wciResponse_9$whas = 1'd1 ;
  assign wci_sfCapSet_9_1$wget = wci_Vm_9_SFlag[0] ;
  assign wci_sfCapSet_9_1$whas = 1'd1 ;
  assign wci_sfCapClear_9_1$wget = 1'd1 ;
  assign wci_sfCapClear_9_1$whas =
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T ;
  assign wci_reqF_10_x_wire$wget = MUX_wci_reqF_10_q_0$write_1__VAL_1 ;
  assign wci_reqF_10_x_wire$whas =
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T ;
  assign wci_wciResponse_10$wget = { wci_Vm_10_SResp, wci_Vm_10_SData } ;
  assign wci_wciResponse_10$whas = 1'd1 ;
  assign wci_sfCapSet_10_1$wget = wci_Vm_10_SFlag[0] ;
  assign wci_sfCapSet_10_1$whas = 1'd1 ;
  assign wci_sfCapClear_10_1$wget = 1'd1 ;
  assign wci_sfCapClear_10_1$whas =
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T ;
  assign wci_reqF_11_x_wire$wget = MUX_wci_reqF_11_q_0$write_1__VAL_1 ;
  assign wci_reqF_11_x_wire$whas =
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T ;
  assign wci_wciResponse_11$wget = { wci_Vm_11_SResp, wci_Vm_11_SData } ;
  assign wci_wciResponse_11$whas = 1'd1 ;
  assign wci_sfCapSet_11_1$wget = wci_Vm_11_SFlag[0] ;
  assign wci_sfCapSet_11_1$whas = 1'd1 ;
  assign wci_sfCapClear_11_1$wget = 1'd1 ;
  assign wci_sfCapClear_11_1$whas =
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T ;
  assign wci_reqF_12_x_wire$wget = MUX_wci_reqF_12_q_0$write_1__VAL_1 ;
  assign wci_reqF_12_x_wire$whas =
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T ;
  assign wci_wciResponse_12$wget = { wci_Vm_12_SResp, wci_Vm_12_SData } ;
  assign wci_wciResponse_12$whas = 1'd1 ;
  assign wci_sfCapSet_12_1$wget = wci_Vm_12_SFlag[0] ;
  assign wci_sfCapSet_12_1$whas = 1'd1 ;
  assign wci_sfCapClear_12_1$wget = 1'd1 ;
  assign wci_sfCapClear_12_1$whas =
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T ;
  assign wci_reqF_13_x_wire$wget = MUX_wci_reqF_13_q_0$write_1__VAL_1 ;
  assign wci_reqF_13_x_wire$whas =
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T ;
  assign wci_wciResponse_13$wget = { wci_Vm_13_SResp, wci_Vm_13_SData } ;
  assign wci_wciResponse_13$whas = 1'd1 ;
  assign wci_sfCapSet_13_1$wget = wci_Vm_13_SFlag[0] ;
  assign wci_sfCapSet_13_1$whas = 1'd1 ;
  assign wci_sfCapClear_13_1$wget = 1'd1 ;
  assign wci_sfCapClear_13_1$whas =
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T ;
  assign wci_reqF_14_x_wire$wget = MUX_wci_reqF_14_q_0$write_1__VAL_1 ;
  assign wci_reqF_14_x_wire$whas =
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T ;
  assign wci_wciResponse_14$wget = { wci_Vm_14_SResp, wci_Vm_14_SData } ;
  assign wci_wciResponse_14$whas = 1'd1 ;
  assign wci_sfCapSet_14_1$wget = wci_Vm_14_SFlag[0] ;
  assign wci_sfCapSet_14_1$whas = 1'd1 ;
  assign wci_sfCapClear_14_1$wget = 1'd1 ;
  assign wci_sfCapClear_14_1$whas =
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T ;
  assign wci_Emv_resp_w$wget = wci_Vm_0_SResp ;
  assign wci_Emv_resp_w$whas = 1'd1 ;
  assign wci_Emv_respData_w$wget = wci_Vm_0_SData ;
  assign wci_Emv_respData_w$whas = 1'd1 ;
  assign wci_Emv_resp_w_1$wget = wci_Vm_1_SResp ;
  assign wci_Emv_resp_w_1$whas = 1'd1 ;
  assign wci_Emv_respData_w_1$wget = wci_Vm_1_SData ;
  assign wci_Emv_respData_w_1$whas = 1'd1 ;
  assign wci_Emv_resp_w_2$wget = wci_Vm_2_SResp ;
  assign wci_Emv_resp_w_2$whas = 1'd1 ;
  assign wci_Emv_respData_w_2$wget = wci_Vm_2_SData ;
  assign wci_Emv_respData_w_2$whas = 1'd1 ;
  assign wci_Emv_resp_w_3$wget = wci_Vm_3_SResp ;
  assign wci_Emv_resp_w_3$whas = 1'd1 ;
  assign wci_Emv_respData_w_3$wget = wci_Vm_3_SData ;
  assign wci_Emv_respData_w_3$whas = 1'd1 ;
  assign wci_Emv_resp_w_4$wget = wci_Vm_4_SResp ;
  assign wci_Emv_resp_w_4$whas = 1'd1 ;
  assign wci_Emv_respData_w_4$wget = wci_Vm_4_SData ;
  assign wci_Emv_respData_w_4$whas = 1'd1 ;
  assign wci_Emv_resp_w_5$wget = wci_Vm_5_SResp ;
  assign wci_Emv_resp_w_5$whas = 1'd1 ;
  assign wci_Emv_respData_w_5$wget = wci_Vm_5_SData ;
  assign wci_Emv_respData_w_5$whas = 1'd1 ;
  assign wci_Emv_resp_w_6$wget = wci_Vm_6_SResp ;
  assign wci_Emv_resp_w_6$whas = 1'd1 ;
  assign wci_Emv_respData_w_6$wget = wci_Vm_6_SData ;
  assign wci_Emv_respData_w_6$whas = 1'd1 ;
  assign wci_Emv_resp_w_7$wget = wci_Vm_7_SResp ;
  assign wci_Emv_resp_w_7$whas = 1'd1 ;
  assign wci_Emv_respData_w_7$wget = wci_Vm_7_SData ;
  assign wci_Emv_respData_w_7$whas = 1'd1 ;
  assign wci_Emv_resp_w_8$wget = wci_Vm_8_SResp ;
  assign wci_Emv_resp_w_8$whas = 1'd1 ;
  assign wci_Emv_respData_w_8$wget = wci_Vm_8_SData ;
  assign wci_Emv_respData_w_8$whas = 1'd1 ;
  assign wci_Emv_resp_w_9$wget = wci_Vm_9_SResp ;
  assign wci_Emv_resp_w_9$whas = 1'd1 ;
  assign wci_Emv_respData_w_9$wget = wci_Vm_9_SData ;
  assign wci_Emv_respData_w_9$whas = 1'd1 ;
  assign wci_Emv_resp_w_10$wget = wci_Vm_10_SResp ;
  assign wci_Emv_resp_w_10$whas = 1'd1 ;
  assign wci_Emv_respData_w_10$wget = wci_Vm_10_SData ;
  assign wci_Emv_respData_w_10$whas = 1'd1 ;
  assign wci_Emv_resp_w_11$wget = wci_Vm_11_SResp ;
  assign wci_Emv_resp_w_11$whas = 1'd1 ;
  assign wci_Emv_respData_w_11$wget = wci_Vm_11_SData ;
  assign wci_Emv_respData_w_11$whas = 1'd1 ;
  assign wci_Emv_resp_w_12$wget = wci_Vm_12_SResp ;
  assign wci_Emv_resp_w_12$whas = 1'd1 ;
  assign wci_Emv_respData_w_12$wget = wci_Vm_12_SData ;
  assign wci_Emv_respData_w_12$whas = 1'd1 ;
  assign wci_Emv_resp_w_13$wget = wci_Vm_13_SResp ;
  assign wci_Emv_resp_w_13$whas = 1'd1 ;
  assign wci_Emv_respData_w_13$wget = wci_Vm_13_SData ;
  assign wci_Emv_respData_w_13$whas = 1'd1 ;
  assign wci_Emv_resp_w_14$wget = wci_Vm_14_SResp ;
  assign wci_Emv_resp_w_14$whas = 1'd1 ;
  assign wci_Emv_respData_w_14$wget = wci_Vm_14_SData ;
  assign wci_Emv_respData_w_14$whas = 1'd1 ;
`ifdef not
  assign rom_serverAdapter_outData_deqCalled$whas =
	     (rom_serverAdapter_outDataCore$EMPTY_N ||
	      rom_serverAdapter_outData_enqData$whas) &&
	     rom_serverAdapter_outData_outData$whas &&
	     adminResp4F$FULL_N ;
`endif
  assign wci_reqF_enqueueing$whas = MUX_wci_busy$write_1__SEL_2 ;
  assign wci_reqF_dequeueing$whas =
	     !wci_sThreadBusy_d && wci_wciResponse$wget[33:32] == 2'd0 &&
	     wci_reqF_c_r ;
  assign wci_sThreadBusy_pw$whas = wci_Vm_0_SThreadBusy ;
  assign wci_reqF_1_enqueueing$whas = MUX_wci_busy_1$write_1__SEL_2 ;
  assign wci_reqF_1_dequeueing$whas =
	     !wci_sThreadBusy_d_1 && wci_wciResponse_1$wget[33:32] == 2'd0 &&
	     wci_reqF_1_c_r ;
  assign wci_sThreadBusy_pw_1$whas = wci_Vm_1_SThreadBusy ;
  assign wci_reqF_2_enqueueing$whas = MUX_wci_busy_2$write_1__SEL_2 ;
  assign wci_reqF_2_dequeueing$whas =
	     !wci_sThreadBusy_d_2 && wci_wciResponse_2$wget[33:32] == 2'd0 &&
	     wci_reqF_2_c_r ;
  assign wci_sThreadBusy_pw_2$whas = wci_Vm_2_SThreadBusy ;
  assign wci_reqF_3_enqueueing$whas = MUX_wci_busy_3$write_1__SEL_2 ;
  assign wci_reqF_3_dequeueing$whas =
	     !wci_sThreadBusy_d_3 && wci_wciResponse_3$wget[33:32] == 2'd0 &&
	     wci_reqF_3_c_r ;
  assign wci_sThreadBusy_pw_3$whas = wci_Vm_3_SThreadBusy ;
  assign wci_reqF_4_enqueueing$whas = MUX_wci_busy_4$write_1__SEL_2 ;
  assign wci_reqF_4_dequeueing$whas =
	     !wci_sThreadBusy_d_4 && wci_wciResponse_4$wget[33:32] == 2'd0 &&
	     wci_reqF_4_c_r ;
  assign wci_sThreadBusy_pw_4$whas = wci_Vm_4_SThreadBusy ;
  assign wci_reqF_5_enqueueing$whas = MUX_wci_busy_5$write_1__SEL_2 ;
  assign wci_reqF_5_dequeueing$whas =
	     !wci_sThreadBusy_d_5 && wci_wciResponse_5$wget[33:32] == 2'd0 &&
	     wci_reqF_5_c_r ;
  assign wci_sThreadBusy_pw_5$whas = wci_Vm_5_SThreadBusy ;
  assign wci_reqF_6_enqueueing$whas = MUX_wci_busy_6$write_1__SEL_2 ;
  assign wci_reqF_6_dequeueing$whas =
	     !wci_sThreadBusy_d_6 && wci_wciResponse_6$wget[33:32] == 2'd0 &&
	     wci_reqF_6_c_r ;
  assign wci_sThreadBusy_pw_6$whas = wci_Vm_6_SThreadBusy ;
  assign wci_reqF_7_enqueueing$whas = MUX_wci_busy_7$write_1__SEL_2 ;
  assign wci_reqF_7_dequeueing$whas =
	     !wci_sThreadBusy_d_7 && wci_wciResponse_7$wget[33:32] == 2'd0 &&
	     wci_reqF_7_c_r ;
  assign wci_sThreadBusy_pw_7$whas = wci_Vm_7_SThreadBusy ;
  assign wci_reqF_8_enqueueing$whas = MUX_wci_busy_8$write_1__SEL_2 ;
  assign wci_reqF_8_dequeueing$whas =
	     !wci_sThreadBusy_d_8 && wci_wciResponse_8$wget[33:32] == 2'd0 &&
	     wci_reqF_8_c_r ;
  assign wci_sThreadBusy_pw_8$whas = wci_Vm_8_SThreadBusy ;
  assign wci_reqF_9_enqueueing$whas = MUX_wci_busy_9$write_1__SEL_2 ;
  assign wci_reqF_9_dequeueing$whas =
	     !wci_sThreadBusy_d_9 && wci_wciResponse_9$wget[33:32] == 2'd0 &&
	     wci_reqF_9_c_r ;
  assign wci_sThreadBusy_pw_9$whas = wci_Vm_9_SThreadBusy ;
  assign wci_reqF_10_enqueueing$whas = MUX_wci_busy_10$write_1__SEL_2 ;
  assign wci_reqF_10_dequeueing$whas =
	     !wci_sThreadBusy_d_10 &&
	     wci_wciResponse_10$wget[33:32] == 2'd0 &&
	     wci_reqF_10_c_r ;
  assign wci_sThreadBusy_pw_10$whas = wci_Vm_10_SThreadBusy ;
  assign wci_reqF_11_enqueueing$whas = MUX_wci_busy_11$write_1__SEL_2 ;
  assign wci_reqF_11_dequeueing$whas =
	     !wci_sThreadBusy_d_11 &&
	     wci_wciResponse_11$wget[33:32] == 2'd0 &&
	     wci_reqF_11_c_r ;
  assign wci_sThreadBusy_pw_11$whas = wci_Vm_11_SThreadBusy ;
  assign wci_reqF_12_enqueueing$whas = MUX_wci_busy_12$write_1__SEL_2 ;
  assign wci_reqF_12_dequeueing$whas =
	     !wci_sThreadBusy_d_12 &&
	     wci_wciResponse_12$wget[33:32] == 2'd0 &&
	     wci_reqF_12_c_r ;
  assign wci_sThreadBusy_pw_12$whas = wci_Vm_12_SThreadBusy ;
  assign wci_reqF_13_enqueueing$whas = MUX_wci_busy_13$write_1__SEL_2 ;
  assign wci_reqF_13_dequeueing$whas =
	     !wci_sThreadBusy_d_13 &&
	     wci_wciResponse_13$wget[33:32] == 2'd0 &&
	     wci_reqF_13_c_r ;
  assign wci_sThreadBusy_pw_13$whas = wci_Vm_13_SThreadBusy ;
  assign wci_reqF_14_enqueueing$whas = MUX_wci_busy_14$write_1__SEL_2 ;
  assign wci_reqF_14_dequeueing$whas =
	     !wci_sThreadBusy_d_14 &&
	     wci_wciResponse_14$wget[33:32] == 2'd0 &&
	     wci_reqF_14_c_r ;
  assign wci_sThreadBusy_pw_14$whas = wci_Vm_14_SThreadBusy ;

  // register cpControl
  assign cpControl$D_IN = cpReq[59:28] ;
  assign cpControl$EN = WILL_FIRE_RL_cpDispatch_T_F_F_T ;

  // register cpReq
  always@(WILL_FIRE_RL_responseAdminRd or
	  WILL_FIRE_RL_cpDispatch_T_F_F_F_F_T_F or
	  WILL_FIRE_RL_cpDispatch_T_F_F_F_F_T_T or
	  WILL_FIRE_RL_reqRcv or
	  MUX_cpReq$write_1__VAL_4 or
	  WILL_FIRE_RL_completeWorkerRead or
	  WILL_FIRE_RL_completeWorkerWrite or
	  WILL_FIRE_RL_cpDispatch_T_F_F_F_F_F_F_F_F_F_F or
	  WILL_FIRE_RL_cpDispatch_T_F_F_F_F_F_F_F_F_F_T or
	  WILL_FIRE_RL_cpDispatch_T_F_F_F_F_F_F_F_F_T or
	  WILL_FIRE_RL_cpDispatch_T_F_F_F_F_F_F_F_T or
	  WILL_FIRE_RL_cpDispatch_T_F_F_F_F_F_F_T or
	  WILL_FIRE_RL_cpDispatch_T_F_F_F_F_F_T or
	  WILL_FIRE_RL_cpDispatch_T_F_F_F_T or
	  WILL_FIRE_RL_cpDispatch_T_F_F_T or
	  WILL_FIRE_RL_cpDispatch_T_F_T or WILL_FIRE_RL_cpDispatch_T_T)
  case (1'b1)
    WILL_FIRE_RL_responseAdminRd || WILL_FIRE_RL_cpDispatch_T_F_F_F_F_T_F ||
    WILL_FIRE_RL_cpDispatch_T_F_F_F_F_T_T:
	cpReq$D_IN = 65'h02AAAAAAAAAAAAAAA;
    WILL_FIRE_RL_reqRcv: cpReq$D_IN = MUX_cpReq$write_1__VAL_4;
    WILL_FIRE_RL_completeWorkerRead || WILL_FIRE_RL_completeWorkerWrite ||
    WILL_FIRE_RL_cpDispatch_T_F_F_F_F_F_F_F_F_F_F ||
    WILL_FIRE_RL_cpDispatch_T_F_F_F_F_F_F_F_F_F_T ||
    WILL_FIRE_RL_cpDispatch_T_F_F_F_F_F_F_F_F_T ||
    WILL_FIRE_RL_cpDispatch_T_F_F_F_F_F_F_F_T ||
    WILL_FIRE_RL_cpDispatch_T_F_F_F_F_F_F_T ||
    WILL_FIRE_RL_cpDispatch_T_F_F_F_F_F_T ||
    WILL_FIRE_RL_cpDispatch_T_F_F_F_T ||
    WILL_FIRE_RL_cpDispatch_T_F_F_T ||
    WILL_FIRE_RL_cpDispatch_T_F_T ||
    WILL_FIRE_RL_cpDispatch_T_T:
	cpReq$D_IN = 65'h02AAAAAAAAAAAAAAA;
    default: cpReq$D_IN = 65'h0AAAAAAAAAAAAAAAA /* unspecified value */ ;
  endcase
  assign cpReq$EN =
	     WILL_FIRE_RL_reqRcv ||
	     WILL_FIRE_RL_cpDispatch_T_F_F_F_F_F_F_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_T_F_F_F_F_F_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_T_F_F_F_F_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_T_F_F_F_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_T_F_F_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_T_F_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_T_F_F_F_F_T_F ||
	     WILL_FIRE_RL_cpDispatch_T_F_F_F_F_T_T ||
	     WILL_FIRE_RL_cpDispatch_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_T_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_T_T ||
	     WILL_FIRE_RL_responseAdminRd ||
	     WILL_FIRE_RL_completeWorkerRead ||
	     WILL_FIRE_RL_completeWorkerWrite ;

  // register deltaTime
`ifdef not
  assign deltaTime$D_IN = timeServ_nowInCC$dD_OUT - { td, cpReq[59:28] } ;
  assign deltaTime$EN = WILL_FIRE_RL_cpDispatch_T_F_F_F_F_F_F_F_F_T ;
`endif

  // register dispatched
  always@(WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_T or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_F or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_F or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_T or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_F or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_F or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_T or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_F or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_F or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_T or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_T_T or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_F or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_F or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_T or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_T_T or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_F or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_F or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_F_T_F_T or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_T_T or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_F_T_F_F or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_F_T_T_F or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_F_T_F_T or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_F_T_T_T or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_T_T or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_F_T_F_F or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_F_T_T_F or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_T_T or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_F_T_F_T or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_F_T_T_T or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_T_T or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_F_T_F_F or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_F_T_T_F or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_F_T_T or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_T_T or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_F_T_F_T or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_F_T_T_T or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_T_T or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_F_T_F_F or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_F_T_T_F or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_F_T_T or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_T_T or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_F_T_F_T or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_F_T_T_T or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_T_T or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_F_T_F_F or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_F_T_T_F or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_F_T_T or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_T_T or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_F_F_T_F_T or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_F_F_T_T_T or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_T_T or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_F_F_T_F_F or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_F_F_T_T_F or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_F_T_T or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_T_T or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_F_F_T_F_T or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_F_F_T_T_T or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_T_T or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_F_F_T_F_F or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_F_F_T_T_F or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_F_T_T or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_T_T or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_F_F_T_F_T or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_F_F_T_T_T or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_T_T or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_F_F_T_F_F or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_F_F_T_T_F or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_F_T_T or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_T_T or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_T_F_F_T_F_T or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_T_F_F_T_T_T or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_T_T_T or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_T_F_F_T_F_F or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_T_F_F_T_T_F or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_T_F_T_T or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_T_T_T or
	  WILL_FIRE_RL_cpDispatch_F_F_T_T_F_F_T_F_T or
	  WILL_FIRE_RL_cpDispatch_F_F_T_T_F_F_T_T_T or
	  WILL_FIRE_RL_cpDispatch_F_F_T_T_T_T or
	  WILL_FIRE_RL_cpDispatch_F_F_T_T_F_F_T_F_F or
	  WILL_FIRE_RL_cpDispatch_F_F_T_T_F_F_T_T_F or
	  WILL_FIRE_RL_cpDispatch_T_F_F_F_F_T_F or
	  WILL_FIRE_RL_cpDispatch_T_F_F_F_F_T_T or
	  WILL_FIRE_RL_reqRcv or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_T_F or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_F_F_T or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_F_T_F or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_T_F or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_F_F_F_T or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_F_F_T or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_F_T_F or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_T_F or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_F_F_F_F_T or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_F_F_F_T or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_F_F_T or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_F_T_F or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_T_F or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_F_F_F_F_F_F or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_F_F_F_F_F_T or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_F_F_F_F_T or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_F_F_F_T or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_F_F_T or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_F_T_F or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_T_F or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_F_F_F_F_F_F or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_F_F_F_F_F_T or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_F_F_F_F_T or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_F_F_F_T or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_F_F_T or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_F_T_F or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_T_F or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_F_F_F_F_F_F or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_F_F_F_F_F_T or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_F_F_F_F_T or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_F_F_F_T or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_F_F_T or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_F_T_F or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_T_F or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_T_F_F_F_F_F_F or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_T_F_F_F_F_F_T or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_T_F_F_F_F_T or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_T_F_F_F_T or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_T_F_F_T or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_T_F_T_F or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_T_T_F or
	  WILL_FIRE_RL_cpDispatch_F_F_F_T or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_T or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_T_F or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_T or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_T_F or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_F_F_F or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_F_F_T or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_T or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_T_F or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_F_F_F or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_F_F_T or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_T or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_T_F or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_F_F_F or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_F_F_T or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_T or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_T_F or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_F_F_F or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_F_F_T or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_T or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_T_F or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_F_F_F or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_F_F_T or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_T or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_T_F or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_F_F_F_F or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_F_F_F_T or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_F_T or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_T_F or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_F_F_F_F or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_F_F_F_T or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_F_T or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_T_F or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_F_F_F_F or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_F_F_F_T or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_F_T or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_T_F or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_T_F_F_F_F or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_T_F_F_F_T or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_T_F_T or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_T_T_F or
	  WILL_FIRE_RL_cpDispatch_F_F_T_T_F_F_F_F or
	  WILL_FIRE_RL_cpDispatch_F_F_T_T_F_F_F_T or
	  WILL_FIRE_RL_cpDispatch_F_F_T_T_F_T or
	  WILL_FIRE_RL_cpDispatch_F_F_T_T_T_F or
`ifdef not
	  WILL_FIRE_RL_rom_serverAdapter_stageReadResponseAlways or
`endif
	  WILL_FIRE_RL_cpDispatch_F_T_F_T or
	  WILL_FIRE_RL_cpDispatch_F_T_T_F_F or
	  WILL_FIRE_RL_cpDispatch_F_T_T_F_T_F_F or
	  WILL_FIRE_RL_cpDispatch_F_T_T_F_T_F_T or
	  WILL_FIRE_RL_cpDispatch_F_T_T_F_T_T or
	  WILL_FIRE_RL_cpDispatch_F_T_T_T or
	  WILL_FIRE_RL_cpDispatch_T_F_F_F_F_F_F_F_F_F_F or
	  WILL_FIRE_RL_cpDispatch_T_F_F_F_F_F_F_F_F_F_T or
	  WILL_FIRE_RL_cpDispatch_T_F_F_F_F_F_F_F_F_T or
	  WILL_FIRE_RL_cpDispatch_T_F_F_F_F_F_F_F_T or
	  WILL_FIRE_RL_cpDispatch_T_F_F_F_F_F_F_T or
	  WILL_FIRE_RL_cpDispatch_T_F_F_F_F_F_T or
	  WILL_FIRE_RL_cpDispatch_T_F_F_F_T or
	  WILL_FIRE_RL_cpDispatch_T_F_F_T or
	  WILL_FIRE_RL_cpDispatch_T_F_T or WILL_FIRE_RL_cpDispatch_T_T)
  case (1'b1)
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_T ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_F ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_F ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_T ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_F ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_F ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_T ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_F ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_F ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_T ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_F ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_F ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_T ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_T_T ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_F ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_F ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_F_T_F_T ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_T_T ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_F_T_F_F ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_F_T_T_F ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_F_T_F_T ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_F_T_T_T ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_T_T ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_F_T_F_F ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_F_T_T_F ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_F_T_F_T ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_F_T_T_T ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_T_T ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_F_T_F_F ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_F_T_T_F ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_F_T_T ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_T_T ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_F_T_F_T ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_F_T_T_T ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_T_T ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_F_T_F_F ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_F_T_T_F ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_F_T_T ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_T_T ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_F_T_F_T ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_F_T_T_T ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_T_T ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_F_T_F_F ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_F_T_T_F ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_F_T_T ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_T_T ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_F_F_T_F_T ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_F_F_T_T_T ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_T_T ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_F_F_T_F_F ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_F_F_T_T_F ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_F_T_T ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_T_T ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_F_F_T_F_T ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_F_F_T_T_T ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_T_T ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_F_F_T_F_F ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_F_F_T_T_F ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_F_T_T ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_T_T ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_F_F_T_F_T ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_F_F_T_T_T ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_T_T ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_F_F_T_F_F ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_F_F_T_T_F ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_F_T_T ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_T_T ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_T_F_F_T_F_T ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_T_F_F_T_T_T ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_T_T_T ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_T_F_F_T_F_F ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_T_F_F_T_T_F ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_T_F_T_T ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_T_T_T ||
    WILL_FIRE_RL_cpDispatch_F_F_T_T_F_F_T_F_T ||
    WILL_FIRE_RL_cpDispatch_F_F_T_T_F_F_T_T_T ||
    WILL_FIRE_RL_cpDispatch_F_F_T_T_T_T ||
    WILL_FIRE_RL_cpDispatch_F_F_T_T_F_F_T_F_F ||
    WILL_FIRE_RL_cpDispatch_F_F_T_T_F_F_T_T_F ||
    WILL_FIRE_RL_cpDispatch_T_F_F_F_F_T_F ||
    WILL_FIRE_RL_cpDispatch_T_F_F_F_F_T_T:
	dispatched$D_IN = 1'd1;
    WILL_FIRE_RL_reqRcv: dispatched$D_IN = 1'd0;
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_T_F ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_F_F_T ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_F_T_F ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_T_F ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_F_F_F_T ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_F_F_T ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_F_T_F ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_T_F ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_F_F_F_F_T ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_F_F_F_T ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_F_F_T ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_F_T_F ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_T_F ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_F_F_F_F_F_F ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_F_F_F_F_F_T ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_F_F_F_F_T ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_F_F_F_T ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_F_F_T ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_F_T_F ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_T_F ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_F_F_F_F_F_F ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_F_F_F_F_F_T ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_F_F_F_F_T ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_F_F_F_T ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_F_F_T ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_F_T_F ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_T_F ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_F_F_F_F_F_F ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_F_F_F_F_F_T ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_F_F_F_F_T ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_F_F_F_T ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_F_F_T ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_F_T_F ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_T_F ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_T_F_F_F_F_F_F ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_T_F_F_F_F_F_T ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_T_F_F_F_F_T ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_T_F_F_F_T ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_T_F_F_T ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_T_F_T_F ||
    WILL_FIRE_RL_cpDispatch_F_F_F_F_T_T_F ||
    WILL_FIRE_RL_cpDispatch_F_F_F_T ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_T ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_T_F ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_T ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_T_F ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_F_F_F ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_F_F_T ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_T ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_T_F ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_F_F_F ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_F_F_T ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_T ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_T_F ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_F_F_F ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_F_F_T ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_T ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_T_F ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_F_F_F ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_F_F_T ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_T ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_T_F ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_F_F_F ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_F_F_T ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_T ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_T_F ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_F_F_F_F ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_F_F_F_T ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_F_T ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_T_F ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_F_F_F_F ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_F_F_F_T ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_F_T ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_T_F ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_F_F_F_F ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_F_F_F_T ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_F_T ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_T_F ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_T_F_F_F_F ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_T_F_F_F_T ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_T_F_T ||
    WILL_FIRE_RL_cpDispatch_F_F_T_F_T_T_F ||
    WILL_FIRE_RL_cpDispatch_F_F_T_T_F_F_F_F ||
    WILL_FIRE_RL_cpDispatch_F_F_T_T_F_F_F_T ||
    WILL_FIRE_RL_cpDispatch_F_F_T_T_F_T ||
    WILL_FIRE_RL_cpDispatch_F_F_T_T_T_F ||
`ifdef not
    WILL_FIRE_RL_rom_serverAdapter_stageReadResponseAlways ||
`endif
    WILL_FIRE_RL_cpDispatch_F_T_F_T ||
    WILL_FIRE_RL_cpDispatch_F_T_T_F_F ||
    WILL_FIRE_RL_cpDispatch_F_T_T_F_T_F_F ||
    WILL_FIRE_RL_cpDispatch_F_T_T_F_T_F_T ||
    WILL_FIRE_RL_cpDispatch_F_T_T_F_T_T ||
    WILL_FIRE_RL_cpDispatch_F_T_T_T ||
    WILL_FIRE_RL_cpDispatch_T_F_F_F_F_F_F_F_F_F_F ||
    WILL_FIRE_RL_cpDispatch_T_F_F_F_F_F_F_F_F_F_T ||
    WILL_FIRE_RL_cpDispatch_T_F_F_F_F_F_F_F_F_T ||
    WILL_FIRE_RL_cpDispatch_T_F_F_F_F_F_F_F_T ||
    WILL_FIRE_RL_cpDispatch_T_F_F_F_F_F_F_T ||
    WILL_FIRE_RL_cpDispatch_T_F_F_F_F_F_T ||
    WILL_FIRE_RL_cpDispatch_T_F_F_F_T ||
    WILL_FIRE_RL_cpDispatch_T_F_F_T ||
    WILL_FIRE_RL_cpDispatch_T_F_T ||
    WILL_FIRE_RL_cpDispatch_T_T:
	dispatched$D_IN = 1'd1;
    default: dispatched$D_IN = 1'b0 /* unspecified value */ ;
  endcase
  assign dispatched$EN =
	     WILL_FIRE_RL_reqRcv ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_F_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_F_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_F_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_F_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_F_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_F_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_F_F_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_F_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_F_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_F_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_F_F_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_F_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_F_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_F_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_F_F_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_F_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_F_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_F_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_T_F_F_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_T_F_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_T_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_T_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_T_F_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_T_F_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_F_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_F_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_F_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_F_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_F_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_F_F_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_F_F_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_F_F_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_T_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_T_F_F_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_T_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_T_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_T_F_F_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_T_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_T_T_T ||
`ifdef not
	     WILL_FIRE_RL_rom_serverAdapter_stageReadResponseAlways ||
`endif
	     WILL_FIRE_RL_cpDispatch_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_T_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_T_T_F_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_T_T_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_T_T_F_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_T_F_F_F_F_F_F_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_T_F_F_F_F_F_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_T_F_F_F_F_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_T_F_F_F_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_T_F_F_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_T_F_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_T_F_F_F_F_T_F ||
	     WILL_FIRE_RL_cpDispatch_T_F_F_F_F_T_T ||
	     WILL_FIRE_RL_cpDispatch_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_T_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_T_T ;

`ifdef not
  // register dna_cnt
  assign dna_cnt$D_IN = dna_cnt + 7'd1 ;
  assign dna_cnt$EN = dna_cnt != 7'd127 ;

  // register dna_rdReg
  assign dna_rdReg$D_IN = dna_rdReg_1$whas ;
  assign dna_rdReg$EN = 1'd1 ;

  // register dna_shftReg
  assign dna_shftReg$D_IN = dna_shftReg_1$whas ;
  assign dna_shftReg$EN = 1'd1 ;

  // register dna_sr
  assign dna_sr$D_IN = { dna_sr[55:0], dna_dna$DOUT } ;
  assign dna_sr$EN = dna_cnt >= 7'd3 && dna_cnt <= 7'd116 && !dna_cnt[0] ;
`endif

  // register readCntReg
  assign readCntReg$D_IN =
	     WILL_FIRE_RL_cpDispatch_T_F_F_F_F_F_F_F_F_F_T ?
	       cpReq[59:28] :
	       MUX_readCntReg$write_1__VAL_2 ;
  assign readCntReg$EN =
	     WILL_FIRE_RL_cpDispatch_T_F_F_F_F_F_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_T_T_F_T_F_T ;

  // register rogueTLP
  assign rogueTLP$D_IN = 4'h0 ;
  assign rogueTLP$EN = 1'b0 ;

`ifdef not
  // register rom_serverAdapter_cnt
  assign rom_serverAdapter_cnt$D_IN =
	     rom_serverAdapter_cnt_29_PLUS_IF_rom_serverAda_ETC___d135 ;
  assign rom_serverAdapter_cnt$EN =
	     WILL_FIRE_RL_rom_serverAdapter_stageReadResponseAlways ||
	     rom_serverAdapter_outData_deqCalled$whas ;

  // register rom_serverAdapter_s1
  assign rom_serverAdapter_s1$D_IN =
	     { WILL_FIRE_RL_rom_serverAdapter_stageReadResponseAlways,
	       1'b1 } ;
  assign rom_serverAdapter_s1$EN = 1'd1 ;
`endif

  // register scratch20
  assign scratch20$D_IN = cpReq[59:28] ;
  assign scratch20$EN = WILL_FIRE_RL_cpDispatch_T_T ;

  // register scratch24
  assign scratch24$D_IN = cpReq[59:28] ;
  assign scratch24$EN = WILL_FIRE_RL_cpDispatch_T_F_T ;

  // register seqTag
  assign seqTag$D_IN = cpReq[35:28] ;
  assign seqTag$EN =
`ifdef not
	     WILL_FIRE_RL_rom_serverAdapter_stageReadResponseAlways ||
`endif
	     WILL_FIRE_RL_cpDispatch_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_T_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_T_T_F_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_T_T_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_T_T_F_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_T_T_T ;

`ifdef not
  // register switch_d
  assign switch_d$D_IN = switch_x ;
  assign switch_d$EN = 1'd1 ;
`endif
  // register td
  assign td$D_IN = cpReq[59:28] ;
  assign td$EN =
	     WILL_FIRE_RL_cpDispatch_T_F_F_F_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_T_F_F_F_F_F_T ;

`ifdef not
  // register timeServ_delSec
  assign timeServ_delSec$D_IN = timeServ_fracSeconds[49:48] ;
  assign timeServ_delSec$EN = 1'd1 ;

  // register timeServ_delSecond
  assign timeServ_delSecond$D_IN =
	     timeServ_fracSeconds - timeServ_lastSecond ;
  assign timeServ_delSecond$EN =
	     timeServ_ppsExtSync_d2 && !timeServ_ppsExtSyncD &&
	     !timeServ_refFromRise_3_ULE_199800000___d5459 &&
	     timeServ_refFromRise_3_ULT_200200000___d5878 ;

  // register timeServ_fracInc
  assign timeServ_fracInc$D_IN = timeServ_fracInc + x__h4421 ;
  assign timeServ_fracInc$EN =
	     timeServ_ppsExtSync_d2_2_AND_NOT_timeServ_ppsE_ETC___d70 ;

  // register timeServ_fracSeconds
  assign timeServ_fracSeconds$D_IN =
	     timeServ_jamFrac ? timeServ_jamFracVal : x__h4649 ;
  assign timeServ_fracSeconds$EN = 1'd1 ;

  // register timeServ_gpsInSticky
  assign timeServ_gpsInSticky$D_IN = 1'd0 ;
  assign timeServ_gpsInSticky$EN = WILL_FIRE_RL_cpDispatch_T_F_F_F_F_T_T ;

  // register timeServ_jamFrac
  assign timeServ_jamFrac$D_IN = timeServ_jamFrac_1$whas ;
  assign timeServ_jamFrac$EN = 1'd1 ;

  // register timeServ_jamFracVal
  assign timeServ_jamFracVal$D_IN =
	     timeServ_jamFrac_1$whas ? x__h3700 : 50'd0 ;
  assign timeServ_jamFracVal$EN = 1'd1 ;

  // register timeServ_lastSecond
  assign timeServ_lastSecond$D_IN = timeServ_fracSeconds ;
  assign timeServ_lastSecond$EN =
	     timeServ_ppsExtSync_d2 && !timeServ_ppsExtSyncD &&
	     !timeServ_refFromRise_3_ULE_199800000___d5459 &&
	     timeServ_refFromRise_3_ULT_200200000___d5878 ;

  // register timeServ_now
  assign timeServ_now$D_IN =
	     { timeServ_refSecCount, timeServ_fracSeconds[47:16] } ;
  assign timeServ_now$EN = timeServ_nowInCC$sRDY ;

  // register timeServ_ppsDrive
  assign timeServ_ppsDrive$D_IN = timeServ_refPerCount < 28'd180000000 ;
  assign timeServ_ppsDrive$EN = 1'd1 ;

  // register timeServ_ppsEdgeCount
  assign timeServ_ppsEdgeCount$D_IN = timeServ_ppsEdgeCount + 8'd1 ;
  assign timeServ_ppsEdgeCount$EN =
	     timeServ_ppsExtSync_d2 && !timeServ_ppsExtSyncD ;

  // register timeServ_ppsExtCapture
  assign timeServ_ppsExtCapture$D_IN = 1'b0 ;
  assign timeServ_ppsExtCapture$EN = 1'b0 ;

  // register timeServ_ppsExtSyncD
  assign timeServ_ppsExtSyncD$D_IN = timeServ_ppsExtSync_d2 ;
  assign timeServ_ppsExtSyncD$EN = !timeServ_ppsDisablePPS$dD_OUT ;

  // register timeServ_ppsExtSync_d1
  assign timeServ_ppsExtSync_d1$D_IN = gps_ppsSyncIn_x ;
  assign timeServ_ppsExtSync_d1$EN = 1'd1 ;

  // register timeServ_ppsExtSync_d2
  assign timeServ_ppsExtSync_d2$D_IN = timeServ_ppsExtSync_d1 ;
  assign timeServ_ppsExtSync_d2$EN = 1'd1 ;

  // register timeServ_ppsInSticky
  assign timeServ_ppsInSticky$D_IN = timeServ_ppsOKCC$dD_OUT ;
  assign timeServ_ppsInSticky$EN =
	     WILL_FIRE_RL_cpDispatch_T_F_F_F_F_T_T ||
	     timeServ_ppsOKCC$dD_OUT ;

  // register timeServ_ppsLost
  assign timeServ_ppsLost$D_IN =
	     timeServ_ppsOK &&
	     timeServ_ppsExtSync_d2_2_AND_NOT_timeServ_ppsE_ETC___d61 ;
  assign timeServ_ppsLost$EN = 1'd1 ;

  // register timeServ_ppsLostSticky
  assign timeServ_ppsLostSticky$D_IN = timeServ_ppsLostCC$dD_OUT ;
  assign timeServ_ppsLostSticky$EN =
	     WILL_FIRE_RL_cpDispatch_T_F_F_F_F_T_T ||
	     timeServ_ppsLostCC$dD_OUT ;

  // register timeServ_ppsOK
  assign timeServ_ppsOK$D_IN =
	     timeServ_ppsExtSync_d2 && !timeServ_ppsExtSyncD &&
	     !timeServ_refFromRise_3_ULE_199800000___d5459 &&
	     timeServ_refFromRise_3_ULT_200200000___d5878 ||
	     timeServ_ppsOK && !timeServ_ppsLost ;
  assign timeServ_ppsOK$EN = 1'd1 ;

  // register timeServ_refFreeCount
  assign timeServ_refFreeCount$D_IN = timeServ_refFreeCount + 28'd1 ;
  assign timeServ_refFreeCount$EN = 1'd1 ;

  // register timeServ_refFreeSamp
  assign timeServ_refFreeSamp$D_IN = timeServ_refFreeCount ;
  assign timeServ_refFreeSamp$EN =
	     timeServ_ppsExtSync_d2 && !timeServ_ppsExtSyncD &&
	     !timeServ_refFromRise_3_ULE_199800000___d5459 &&
	     timeServ_refFromRise_3_ULT_200200000___d5878 ;

  // register timeServ_refFreeSpan
  assign timeServ_refFreeSpan$D_IN =
	     timeServ_refFreeCount - timeServ_refFreeSamp ;
  assign timeServ_refFreeSpan$EN =
	     timeServ_ppsExtSync_d2 && !timeServ_ppsExtSyncD &&
	     !timeServ_refFromRise_3_ULE_199800000___d5459 &&
	     timeServ_refFromRise_3_ULT_200200000___d5878 ;

  // register timeServ_refFromRise
  assign timeServ_refFromRise$D_IN =
	     (timeServ_ppsExtSync_d2 && !timeServ_ppsExtSyncD) ?
	       28'd0 :
	       timeServ_refFromRise + 28'd1 ;
  assign timeServ_refFromRise$EN = 1'd1 ;

  // register timeServ_refPerCount
  assign timeServ_refPerCount$D_IN =
	     IF_timeServ_ppsOK_7_THEN_timeServ_ppsExtSync_d_ETC___d5465 ?
	       28'd0 :
	       timeServ_refPerCount + 28'd1 ;
  assign timeServ_refPerCount$EN = 1'd1 ;

  // register timeServ_refSecCount
  assign timeServ_refSecCount$D_IN =
	     timeServ_setRefF$dEMPTY_N ?
	       timeServ_setRefF$dD_OUT[63:32] :
	       x__h4715 ;
  assign timeServ_refSecCount$EN =
	     timeServ_setRefF$dEMPTY_N ||
	     IF_timeServ_ppsOK_7_THEN_timeServ_ppsExtSync_d_ETC___d5465 ;

  // register timeServ_rplTimeControl
  assign timeServ_rplTimeControl$D_IN = cpReq[32:28] ;
  assign timeServ_rplTimeControl$EN =
	     WILL_FIRE_RL_cpDispatch_T_F_F_F_F_T_F ||
	     WILL_FIRE_RL_cpDispatch_T_F_F_F_F_T_T ;

  // register timeServ_timeSetSticky
  assign timeServ_timeSetSticky$D_IN =
	     !WILL_FIRE_RL_cpDispatch_T_F_F_F_F_T_T ;
  assign timeServ_timeSetSticky$EN =
	     WILL_FIRE_RL_cpDispatch_T_F_F_F_F_T_T ||
	     WILL_FIRE_RL_cpDispatch_T_F_F_F_F_F_F_T ;

  // register timeServ_xo2
  assign timeServ_xo2$D_IN = !timeServ_xo2 ;
  assign timeServ_xo2$EN = 1'd1 ;
`endif

  // register warmResetP
  assign warmResetP$D_IN =
	     WILL_FIRE_RL_cpDispatch_T_F_F_F_T &&
	     cpReq[59:28] == 32'hC0DEFFFF ;
  assign warmResetP$EN = 1'd1 ;

  // register wci_busy
  assign wci_busy$D_IN = !MUX_wci_busy$write_1__SEL_1 ;
  assign wci_busy$EN =
	     WILL_FIRE_RL_wci_wrkBusy &&
	     (!wci_respTimr_28_ULT_1_SL_wci_wTimeout_29_30___d5879 ||
	      wci_wciResponse$wget[33:32] != 2'd0) ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_T_F_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_T_T_T ;

  // register wci_busy_1
  assign wci_busy_1$D_IN = !MUX_wci_busy_1$write_1__SEL_1 ;
  assign wci_busy_1$EN =
	     WILL_FIRE_RL_wci_wrkBusy_1 &&
	     (!wci_respTimr_1_68_ULT_1_SL_wci_wTimeout_1_69_70___d5880 ||
	      wci_wciResponse_1$wget[33:32] != 2'd0) ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_F_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_T_T_T ;

  // register wci_busy_10
  assign wci_busy_10$D_IN = !MUX_wci_busy_10$write_1__SEL_1 ;
  assign wci_busy_10$EN =
	     WILL_FIRE_RL_wci_wrkBusy_10 &&
	     (!wci_respTimr_10_628_ULT_1_SL_wci_wTimeout_10_6_ETC___d5889 ||
	      wci_wciResponse_10$wget[33:32] != 2'd0) ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_T_T ;

  // register wci_busy_11
  assign wci_busy_11$D_IN = !MUX_wci_busy_11$write_1__SEL_1 ;
  assign wci_busy_11$EN =
	     WILL_FIRE_RL_wci_wrkBusy_11 &&
	     (!wci_respTimr_11_768_ULT_1_SL_wci_wTimeout_11_7_ETC___d5890 ||
	      wci_wciResponse_11$wget[33:32] != 2'd0) ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_T_T ;

  // register wci_busy_12
  assign wci_busy_12$D_IN = !MUX_wci_busy_12$write_1__SEL_1 ;
  assign wci_busy_12$EN =
	     WILL_FIRE_RL_wci_wrkBusy_12 &&
	     (!wci_respTimr_12_908_ULT_1_SL_wci_wTimeout_12_9_ETC___d5891 ||
	      wci_wciResponse_12$wget[33:32] != 2'd0) ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ;

  // register wci_busy_13
  assign wci_busy_13$D_IN = !MUX_wci_busy_13$write_1__SEL_1 ;
  assign wci_busy_13$EN =
	     WILL_FIRE_RL_wci_wrkBusy_13 &&
	     (!wci_respTimr_13_048_ULT_1_SL_wci_wTimeout_13_0_ETC___d5892 ||
	      wci_wciResponse_13$wget[33:32] != 2'd0) ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ;

  // register wci_busy_14
  assign wci_busy_14$D_IN = !MUX_wci_busy_14$write_1__SEL_1 ;
  assign wci_busy_14$EN =
	     WILL_FIRE_RL_wci_wrkBusy_14 &&
	     (!wci_respTimr_14_188_ULT_1_SL_wci_wTimeout_14_1_ETC___d5893 ||
	      wci_wciResponse_14$wget[33:32] != 2'd0) ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ;

  // register wci_busy_2
  assign wci_busy_2$D_IN = !MUX_wci_busy_2$write_1__SEL_1 ;
  assign wci_busy_2$EN =
	     WILL_FIRE_RL_wci_wrkBusy_2 &&
	     (!wci_respTimr_2_08_ULT_1_SL_wci_wTimeout_2_09_10___d5881 ||
	      wci_wciResponse_2$wget[33:32] != 2'd0) ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_F_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_T_T ;

  // register wci_busy_3
  assign wci_busy_3$D_IN = !MUX_wci_busy_3$write_1__SEL_1 ;
  assign wci_busy_3$EN =
	     WILL_FIRE_RL_wci_wrkBusy_3 &&
	     (!wci_respTimr_3_48_ULT_1_SL_wci_wTimeout_3_49_50___d5882 ||
	      wci_wciResponse_3$wget[33:32] != 2'd0) ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_F_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_T_T ;

  // register wci_busy_4
  assign wci_busy_4$D_IN = !MUX_wci_busy_4$write_1__SEL_1 ;
  assign wci_busy_4$EN =
	     WILL_FIRE_RL_wci_wrkBusy_4 &&
	     (!wci_respTimr_4_88_ULT_1_SL_wci_wTimeout_4_89_90___d5883 ||
	      wci_wciResponse_4$wget[33:32] != 2'd0) ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_F_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_T_T ;

  // register wci_busy_5
  assign wci_busy_5$D_IN = !MUX_wci_busy_5$write_1__SEL_1 ;
  assign wci_busy_5$EN =
	     WILL_FIRE_RL_wci_wrkBusy_5 &&
	     (!wci_respTimr_5_28_ULT_1_SL_wci_wTimeout_5_29_30___d5884 ||
	      wci_wciResponse_5$wget[33:32] != 2'd0) ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_F_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_T_T ;

  // register wci_busy_6
  assign wci_busy_6$D_IN = !MUX_wci_busy_6$write_1__SEL_1 ;
  assign wci_busy_6$EN =
	     WILL_FIRE_RL_wci_wrkBusy_6 &&
	     (!wci_respTimr_6_068_ULT_1_SL_wci_wTimeout_6_069_ETC___d5885 ||
	      wci_wciResponse_6$wget[33:32] != 2'd0) ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_F_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_T_T ;

  // register wci_busy_7
  assign wci_busy_7$D_IN = !MUX_wci_busy_7$write_1__SEL_1 ;
  assign wci_busy_7$EN =
	     WILL_FIRE_RL_wci_wrkBusy_7 &&
	     (!wci_respTimr_7_208_ULT_1_SL_wci_wTimeout_7_209_ETC___d5886 ||
	      wci_wciResponse_7$wget[33:32] != 2'd0) ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_T_T ;

  // register wci_busy_8
  assign wci_busy_8$D_IN = !MUX_wci_busy_8$write_1__SEL_1 ;
  assign wci_busy_8$EN =
	     WILL_FIRE_RL_wci_wrkBusy_8 &&
	     (!wci_respTimr_8_348_ULT_1_SL_wci_wTimeout_8_349_ETC___d5887 ||
	      wci_wciResponse_8$wget[33:32] != 2'd0) ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_T_T ;

  // register wci_busy_9
  assign wci_busy_9$D_IN = !MUX_wci_busy_9$write_1__SEL_1 ;
  assign wci_busy_9$EN =
	     WILL_FIRE_RL_wci_wrkBusy_9 &&
	     (!wci_respTimr_9_488_ULT_1_SL_wci_wTimeout_9_489_ETC___d5888 ||
	      wci_wciResponse_9$wget[33:32] != 2'd0) ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_T_T ;

  // register wci_lastConfigAddr
  assign wci_lastConfigAddr$D_IN = { 13'd4096, cpReq[23:4] } ;
  assign wci_lastConfigAddr$EN =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_T_T_T ;

  // register wci_lastConfigAddr_1
  assign wci_lastConfigAddr_1$D_IN = wci_lastConfigAddr$D_IN ;
  assign wci_lastConfigAddr_1$EN =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_T_T_T ;

  // register wci_lastConfigAddr_10
  assign wci_lastConfigAddr_10$D_IN = wci_lastConfigAddr$D_IN ;
  assign wci_lastConfigAddr_10$EN =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_T_T ;

  // register wci_lastConfigAddr_11
  assign wci_lastConfigAddr_11$D_IN = wci_lastConfigAddr$D_IN ;
  assign wci_lastConfigAddr_11$EN =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_T_T ;

  // register wci_lastConfigAddr_12
  assign wci_lastConfigAddr_12$D_IN = wci_lastConfigAddr$D_IN ;
  assign wci_lastConfigAddr_12$EN =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ;

  // register wci_lastConfigAddr_13
  assign wci_lastConfigAddr_13$D_IN = wci_lastConfigAddr$D_IN ;
  assign wci_lastConfigAddr_13$EN =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ;

  // register wci_lastConfigAddr_14
  assign wci_lastConfigAddr_14$D_IN = wci_lastConfigAddr$D_IN ;
  assign wci_lastConfigAddr_14$EN =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ;

  // register wci_lastConfigAddr_2
  assign wci_lastConfigAddr_2$D_IN = wci_lastConfigAddr$D_IN ;
  assign wci_lastConfigAddr_2$EN =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_T_T ;

  // register wci_lastConfigAddr_3
  assign wci_lastConfigAddr_3$D_IN = wci_lastConfigAddr$D_IN ;
  assign wci_lastConfigAddr_3$EN =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_T_T ;

  // register wci_lastConfigAddr_4
  assign wci_lastConfigAddr_4$D_IN = wci_lastConfigAddr$D_IN ;
  assign wci_lastConfigAddr_4$EN =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_T_T ;

  // register wci_lastConfigAddr_5
  assign wci_lastConfigAddr_5$D_IN = wci_lastConfigAddr$D_IN ;
  assign wci_lastConfigAddr_5$EN =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_T_T ;

  // register wci_lastConfigAddr_6
  assign wci_lastConfigAddr_6$D_IN = wci_lastConfigAddr$D_IN ;
  assign wci_lastConfigAddr_6$EN =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_T_T ;

  // register wci_lastConfigAddr_7
  assign wci_lastConfigAddr_7$D_IN = wci_lastConfigAddr$D_IN ;
  assign wci_lastConfigAddr_7$EN =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_T_T ;

  // register wci_lastConfigAddr_8
  assign wci_lastConfigAddr_8$D_IN = wci_lastConfigAddr$D_IN ;
  assign wci_lastConfigAddr_8$EN =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_T_T ;

  // register wci_lastConfigAddr_9
  assign wci_lastConfigAddr_9$D_IN = wci_lastConfigAddr$D_IN ;
  assign wci_lastConfigAddr_9$EN =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_T_T ;

  // register wci_lastConfigBE
  assign wci_lastConfigBE$D_IN = { 1'd1, cpReq[3:0] } ;
  assign wci_lastConfigBE$EN =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_T_T_T ;

  // register wci_lastConfigBE_1
  assign wci_lastConfigBE_1$D_IN = wci_lastConfigBE$D_IN ;
  assign wci_lastConfigBE_1$EN =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_T_T_T ;

  // register wci_lastConfigBE_10
  assign wci_lastConfigBE_10$D_IN = wci_lastConfigBE$D_IN ;
  assign wci_lastConfigBE_10$EN =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_T_T ;

  // register wci_lastConfigBE_11
  assign wci_lastConfigBE_11$D_IN = wci_lastConfigBE$D_IN ;
  assign wci_lastConfigBE_11$EN =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_T_T ;

  // register wci_lastConfigBE_12
  assign wci_lastConfigBE_12$D_IN = wci_lastConfigBE$D_IN ;
  assign wci_lastConfigBE_12$EN =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ;

  // register wci_lastConfigBE_13
  assign wci_lastConfigBE_13$D_IN = wci_lastConfigBE$D_IN ;
  assign wci_lastConfigBE_13$EN =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ;

  // register wci_lastConfigBE_14
  assign wci_lastConfigBE_14$D_IN = wci_lastConfigBE$D_IN ;
  assign wci_lastConfigBE_14$EN =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ;

  // register wci_lastConfigBE_2
  assign wci_lastConfigBE_2$D_IN = wci_lastConfigBE$D_IN ;
  assign wci_lastConfigBE_2$EN =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_T_T ;

  // register wci_lastConfigBE_3
  assign wci_lastConfigBE_3$D_IN = wci_lastConfigBE$D_IN ;
  assign wci_lastConfigBE_3$EN =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_T_T ;

  // register wci_lastConfigBE_4
  assign wci_lastConfigBE_4$D_IN = wci_lastConfigBE$D_IN ;
  assign wci_lastConfigBE_4$EN =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_T_T ;

  // register wci_lastConfigBE_5
  assign wci_lastConfigBE_5$D_IN = wci_lastConfigBE$D_IN ;
  assign wci_lastConfigBE_5$EN =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_T_T ;

  // register wci_lastConfigBE_6
  assign wci_lastConfigBE_6$D_IN = wci_lastConfigBE$D_IN ;
  assign wci_lastConfigBE_6$EN =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_T_T ;

  // register wci_lastConfigBE_7
  assign wci_lastConfigBE_7$D_IN = wci_lastConfigBE$D_IN ;
  assign wci_lastConfigBE_7$EN =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_T_T ;

  // register wci_lastConfigBE_8
  assign wci_lastConfigBE_8$D_IN = wci_lastConfigBE$D_IN ;
  assign wci_lastConfigBE_8$EN =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_T_T ;

  // register wci_lastConfigBE_9
  assign wci_lastConfigBE_9$D_IN = wci_lastConfigBE$D_IN ;
  assign wci_lastConfigBE_9$EN =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_T_T ;

  // register wci_lastControlOp
  assign wci_lastControlOp$D_IN = { 1'd1, cpReq[8:6] } ;
  assign wci_lastControlOp$EN = WILL_FIRE_RL_cpDispatch_F_F_F_F_T_F_T_T ;

  // register wci_lastControlOp_1
  assign wci_lastControlOp_1$D_IN = wci_lastControlOp$D_IN ;
  assign wci_lastControlOp_1$EN = WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_F_T_T ;

  // register wci_lastControlOp_10
  assign wci_lastControlOp_10$D_IN = wci_lastControlOp$D_IN ;
  assign wci_lastControlOp_10$EN =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T ;

  // register wci_lastControlOp_11
  assign wci_lastControlOp_11$D_IN = wci_lastControlOp$D_IN ;
  assign wci_lastControlOp_11$EN =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T ;

  // register wci_lastControlOp_12
  assign wci_lastControlOp_12$D_IN = wci_lastControlOp$D_IN ;
  assign wci_lastControlOp_12$EN =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T ;

  // register wci_lastControlOp_13
  assign wci_lastControlOp_13$D_IN = wci_lastControlOp$D_IN ;
  assign wci_lastControlOp_13$EN =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T ;

  // register wci_lastControlOp_14
  assign wci_lastControlOp_14$D_IN = wci_lastControlOp$D_IN ;
  assign wci_lastControlOp_14$EN =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T ;

  // register wci_lastControlOp_2
  assign wci_lastControlOp_2$D_IN = wci_lastControlOp$D_IN ;
  assign wci_lastControlOp_2$EN =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_F_T_T ;

  // register wci_lastControlOp_3
  assign wci_lastControlOp_3$D_IN = wci_lastControlOp$D_IN ;
  assign wci_lastControlOp_3$EN =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_F_T_T ;

  // register wci_lastControlOp_4
  assign wci_lastControlOp_4$D_IN = wci_lastControlOp$D_IN ;
  assign wci_lastControlOp_4$EN =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_F_T_T ;

  // register wci_lastControlOp_5
  assign wci_lastControlOp_5$D_IN = wci_lastControlOp$D_IN ;
  assign wci_lastControlOp_5$EN =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_F_T_T ;

  // register wci_lastControlOp_6
  assign wci_lastControlOp_6$D_IN = wci_lastControlOp$D_IN ;
  assign wci_lastControlOp_6$EN =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_F_T_T ;

  // register wci_lastControlOp_7
  assign wci_lastControlOp_7$D_IN = wci_lastControlOp$D_IN ;
  assign wci_lastControlOp_7$EN =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T ;

  // register wci_lastControlOp_8
  assign wci_lastControlOp_8$D_IN = wci_lastControlOp$D_IN ;
  assign wci_lastControlOp_8$EN =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T ;

  // register wci_lastControlOp_9
  assign wci_lastControlOp_9$D_IN = wci_lastControlOp$D_IN ;
  assign wci_lastControlOp_9$EN =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T ;

  // register wci_lastOpWrite
  assign wci_lastOpWrite$D_IN =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_T_T_T ? 2'd2 : 2'd3 ;
  assign wci_lastOpWrite$EN =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_T_T_T ;

  // register wci_lastOpWrite_1
  assign wci_lastOpWrite_1$D_IN =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_T_T ? 2'd2 : 2'd3 ;
  assign wci_lastOpWrite_1$EN =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_T_T_T ;

  // register wci_lastOpWrite_10
  assign wci_lastOpWrite_10$D_IN =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ?
	       2'd2 :
	       2'd3 ;
  assign wci_lastOpWrite_10$EN =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_T_T ;

  // register wci_lastOpWrite_11
  assign wci_lastOpWrite_11$D_IN =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ?
	       2'd2 :
	       2'd3 ;
  assign wci_lastOpWrite_11$EN =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_T_T ;

  // register wci_lastOpWrite_12
  assign wci_lastOpWrite_12$D_IN =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ?
	       2'd2 :
	       2'd3 ;
  assign wci_lastOpWrite_12$EN =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ;

  // register wci_lastOpWrite_13
  assign wci_lastOpWrite_13$D_IN =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ?
	       2'd2 :
	       2'd3 ;
  assign wci_lastOpWrite_13$EN =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ;

  // register wci_lastOpWrite_14
  assign wci_lastOpWrite_14$D_IN =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ?
	       2'd2 :
	       2'd3 ;
  assign wci_lastOpWrite_14$EN =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ;

  // register wci_lastOpWrite_2
  assign wci_lastOpWrite_2$D_IN =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_T_T ? 2'd2 : 2'd3 ;
  assign wci_lastOpWrite_2$EN =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_T_T ;

  // register wci_lastOpWrite_3
  assign wci_lastOpWrite_3$D_IN =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_T_T ? 2'd2 : 2'd3 ;
  assign wci_lastOpWrite_3$EN =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_T_T ;

  // register wci_lastOpWrite_4
  assign wci_lastOpWrite_4$D_IN =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_T_T ? 2'd2 : 2'd3 ;
  assign wci_lastOpWrite_4$EN =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_T_T ;

  // register wci_lastOpWrite_5
  assign wci_lastOpWrite_5$D_IN =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_T_T ? 2'd2 : 2'd3 ;
  assign wci_lastOpWrite_5$EN =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_T_T ;

  // register wci_lastOpWrite_6
  assign wci_lastOpWrite_6$D_IN =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_T_T ? 2'd2 : 2'd3 ;
  assign wci_lastOpWrite_6$EN =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_T_T ;

  // register wci_lastOpWrite_7
  assign wci_lastOpWrite_7$D_IN =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_T_T ?
	       2'd2 :
	       2'd3 ;
  assign wci_lastOpWrite_7$EN =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_T_T ;

  // register wci_lastOpWrite_8
  assign wci_lastOpWrite_8$D_IN =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ?
	       2'd2 :
	       2'd3 ;
  assign wci_lastOpWrite_8$EN =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_T_T ;

  // register wci_lastOpWrite_9
  assign wci_lastOpWrite_9$D_IN =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ?
	       2'd2 :
	       2'd3 ;
  assign wci_lastOpWrite_9$EN =
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_T_T ;

  // register wci_mFlagReg
  assign wci_mFlagReg$D_IN = 2'h0 ;
  assign wci_mFlagReg$EN = 1'b0 ;

  // register wci_mFlagReg_1
  assign wci_mFlagReg_1$D_IN = 2'h0 ;
  assign wci_mFlagReg_1$EN = 1'b0 ;

  // register wci_mFlagReg_10
  assign wci_mFlagReg_10$D_IN = 2'h0 ;
  assign wci_mFlagReg_10$EN = 1'b0 ;

  // register wci_mFlagReg_11
  assign wci_mFlagReg_11$D_IN = 2'h0 ;
  assign wci_mFlagReg_11$EN = 1'b0 ;

  // register wci_mFlagReg_12
  assign wci_mFlagReg_12$D_IN = 2'h0 ;
  assign wci_mFlagReg_12$EN = 1'b0 ;

  // register wci_mFlagReg_13
  assign wci_mFlagReg_13$D_IN = 2'h0 ;
  assign wci_mFlagReg_13$EN = 1'b0 ;

  // register wci_mFlagReg_14
  assign wci_mFlagReg_14$D_IN = 2'h0 ;
  assign wci_mFlagReg_14$EN = 1'b0 ;

  // register wci_mFlagReg_2
  assign wci_mFlagReg_2$D_IN = 2'h0 ;
  assign wci_mFlagReg_2$EN = 1'b0 ;

  // register wci_mFlagReg_3
  assign wci_mFlagReg_3$D_IN = 2'h0 ;
  assign wci_mFlagReg_3$EN = 1'b0 ;

  // register wci_mFlagReg_4
  assign wci_mFlagReg_4$D_IN = 2'h0 ;
  assign wci_mFlagReg_4$EN = 1'b0 ;

  // register wci_mFlagReg_5
  assign wci_mFlagReg_5$D_IN = 2'h0 ;
  assign wci_mFlagReg_5$EN = 1'b0 ;

  // register wci_mFlagReg_6
  assign wci_mFlagReg_6$D_IN = 2'h0 ;
  assign wci_mFlagReg_6$EN = 1'b0 ;

  // register wci_mFlagReg_7
  assign wci_mFlagReg_7$D_IN = 2'h0 ;
  assign wci_mFlagReg_7$EN = 1'b0 ;

  // register wci_mFlagReg_8
  assign wci_mFlagReg_8$D_IN = 2'h0 ;
  assign wci_mFlagReg_8$EN = 1'b0 ;

  // register wci_mFlagReg_9
  assign wci_mFlagReg_9$D_IN = 2'h0 ;
  assign wci_mFlagReg_9$EN = 1'b0 ;

  // register wci_pageWindow
  assign wci_pageWindow$D_IN = cpReq[39:28] ;
  assign wci_pageWindow$EN = WILL_FIRE_RL_cpDispatch_F_F_T_T_F_F_F_T ;

  // register wci_pageWindow_1
  assign wci_pageWindow_1$D_IN = cpReq[39:28] ;
  assign wci_pageWindow_1$EN = WILL_FIRE_RL_cpDispatch_F_F_T_F_T_F_F_F_T ;

  // register wci_pageWindow_10
  assign wci_pageWindow_10$D_IN = cpReq[39:28] ;
  assign wci_pageWindow_10$EN =
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T ;

  // register wci_pageWindow_11
  assign wci_pageWindow_11$D_IN = cpReq[39:28] ;
  assign wci_pageWindow_11$EN =
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T ;

  // register wci_pageWindow_12
  assign wci_pageWindow_12$D_IN = cpReq[39:28] ;
  assign wci_pageWindow_12$EN =
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T ;

  // register wci_pageWindow_13
  assign wci_pageWindow_13$D_IN = cpReq[39:28] ;
  assign wci_pageWindow_13$EN =
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T ;

  // register wci_pageWindow_14
  assign wci_pageWindow_14$D_IN = cpReq[39:28] ;
  assign wci_pageWindow_14$EN =
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T ;

  // register wci_pageWindow_2
  assign wci_pageWindow_2$D_IN = cpReq[39:28] ;
  assign wci_pageWindow_2$EN = WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_F_F_F_T ;

  // register wci_pageWindow_3
  assign wci_pageWindow_3$D_IN = cpReq[39:28] ;
  assign wci_pageWindow_3$EN = WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_F_F_F_T ;

  // register wci_pageWindow_4
  assign wci_pageWindow_4$D_IN = cpReq[39:28] ;
  assign wci_pageWindow_4$EN =
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_F_F_F_T ;

  // register wci_pageWindow_5
  assign wci_pageWindow_5$D_IN = cpReq[39:28] ;
  assign wci_pageWindow_5$EN =
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_F_F_T ;

  // register wci_pageWindow_6
  assign wci_pageWindow_6$D_IN = cpReq[39:28] ;
  assign wci_pageWindow_6$EN =
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_F_F_T ;

  // register wci_pageWindow_7
  assign wci_pageWindow_7$D_IN = cpReq[39:28] ;
  assign wci_pageWindow_7$EN =
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_F_F_T ;

  // register wci_pageWindow_8
  assign wci_pageWindow_8$D_IN = cpReq[39:28] ;
  assign wci_pageWindow_8$EN =
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_F_F_T ;

  // register wci_pageWindow_9
  assign wci_pageWindow_9$D_IN = cpReq[39:28] ;
  assign wci_pageWindow_9$EN =
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_F_F_T ;

  // register wci_reqERR
  assign wci_reqERR$D_IN =
	     MUX_wci_reqERR$write_1__SEL_1 ?
	       MUX_wci_reqERR$write_1__VAL_1 :
	       3'd0 ;
  assign wci_reqERR$EN =
	     WILL_FIRE_RL_wci_wrkBusy &&
	     wci_wciResponse$wget[33:32] == 2'd3 &&
	     (wci_reqPend == 2'd1 || wci_reqPend == 2'd2 ||
	      wci_reqPend == 2'd3) ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_T_F_F_T_T_T ;

  // register wci_reqERR_1
  assign wci_reqERR_1$D_IN =
	     MUX_wci_reqERR_1$write_1__SEL_1 ?
	       MUX_wci_reqERR_1$write_1__VAL_1 :
	       3'd0 ;
  assign wci_reqERR_1$EN =
	     WILL_FIRE_RL_wci_wrkBusy_1 &&
	     wci_wciResponse_1$wget[33:32] == 2'd3 &&
	     (wci_reqPend_1 == 2'd1 || wci_reqPend_1 == 2'd2 ||
	      wci_reqPend_1 == 2'd3) ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_T_F_F_T_T_T ;

  // register wci_reqERR_10
  assign wci_reqERR_10$D_IN =
	     MUX_wci_reqERR_10$write_1__SEL_1 ?
	       MUX_wci_reqERR_10$write_1__VAL_1 :
	       3'd0 ;
  assign wci_reqERR_10$EN =
	     WILL_FIRE_RL_wci_wrkBusy_10 &&
	     wci_wciResponse_10$wget[33:32] == 2'd3 &&
	     (wci_reqPend_10 == 2'd1 || wci_reqPend_10 == 2'd2 ||
	      wci_reqPend_10 == 2'd3) ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T ;

  // register wci_reqERR_11
  assign wci_reqERR_11$D_IN =
	     MUX_wci_reqERR_11$write_1__SEL_1 ?
	       MUX_wci_reqERR_11$write_1__VAL_1 :
	       3'd0 ;
  assign wci_reqERR_11$EN =
	     WILL_FIRE_RL_wci_wrkBusy_11 &&
	     wci_wciResponse_11$wget[33:32] == 2'd3 &&
	     (wci_reqPend_11 == 2'd1 || wci_reqPend_11 == 2'd2 ||
	      wci_reqPend_11 == 2'd3) ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T ;

  // register wci_reqERR_12
  assign wci_reqERR_12$D_IN =
	     MUX_wci_reqERR_12$write_1__SEL_1 ?
	       MUX_wci_reqERR_12$write_1__VAL_1 :
	       3'd0 ;
  assign wci_reqERR_12$EN =
	     WILL_FIRE_RL_wci_wrkBusy_12 &&
	     wci_wciResponse_12$wget[33:32] == 2'd3 &&
	     (wci_reqPend_12 == 2'd1 || wci_reqPend_12 == 2'd2 ||
	      wci_reqPend_12 == 2'd3) ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T ;

  // register wci_reqERR_13
  assign wci_reqERR_13$D_IN =
	     MUX_wci_reqERR_13$write_1__SEL_1 ?
	       MUX_wci_reqERR_13$write_1__VAL_1 :
	       3'd0 ;
  assign wci_reqERR_13$EN =
	     WILL_FIRE_RL_wci_wrkBusy_13 &&
	     wci_wciResponse_13$wget[33:32] == 2'd3 &&
	     (wci_reqPend_13 == 2'd1 || wci_reqPend_13 == 2'd2 ||
	      wci_reqPend_13 == 2'd3) ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T ;

  // register wci_reqERR_14
  assign wci_reqERR_14$D_IN =
	     MUX_wci_reqERR_14$write_1__SEL_1 ?
	       MUX_wci_reqERR_14$write_1__VAL_1 :
	       3'd0 ;
  assign wci_reqERR_14$EN =
	     WILL_FIRE_RL_wci_wrkBusy_14 &&
	     wci_wciResponse_14$wget[33:32] == 2'd3 &&
	     (wci_reqPend_14 == 2'd1 || wci_reqPend_14 == 2'd2 ||
	      wci_reqPend_14 == 2'd3) ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T ;

  // register wci_reqERR_2
  assign wci_reqERR_2$D_IN =
	     MUX_wci_reqERR_2$write_1__SEL_1 ?
	       MUX_wci_reqERR_2$write_1__VAL_1 :
	       3'd0 ;
  assign wci_reqERR_2$EN =
	     WILL_FIRE_RL_wci_wrkBusy_2 &&
	     wci_wciResponse_2$wget[33:32] == 2'd3 &&
	     (wci_reqPend_2 == 2'd1 || wci_reqPend_2 == 2'd2 ||
	      wci_reqPend_2 == 2'd3) ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_F_F_T_T_T ;

  // register wci_reqERR_3
  assign wci_reqERR_3$D_IN =
	     MUX_wci_reqERR_3$write_1__SEL_1 ?
	       MUX_wci_reqERR_3$write_1__VAL_1 :
	       3'd0 ;
  assign wci_reqERR_3$EN =
	     WILL_FIRE_RL_wci_wrkBusy_3 &&
	     wci_wciResponse_3$wget[33:32] == 2'd3 &&
	     (wci_reqPend_3 == 2'd1 || wci_reqPend_3 == 2'd2 ||
	      wci_reqPend_3 == 2'd3) ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_F_F_T_T_T ;

  // register wci_reqERR_4
  assign wci_reqERR_4$D_IN =
	     MUX_wci_reqERR_4$write_1__SEL_1 ?
	       MUX_wci_reqERR_4$write_1__VAL_1 :
	       3'd0 ;
  assign wci_reqERR_4$EN =
	     WILL_FIRE_RL_wci_wrkBusy_4 &&
	     wci_wciResponse_4$wget[33:32] == 2'd3 &&
	     (wci_reqPend_4 == 2'd1 || wci_reqPend_4 == 2'd2 ||
	      wci_reqPend_4 == 2'd3) ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_F_F_T_T_T ;

  // register wci_reqERR_5
  assign wci_reqERR_5$D_IN =
	     MUX_wci_reqERR_5$write_1__SEL_1 ?
	       MUX_wci_reqERR_5$write_1__VAL_1 :
	       3'd0 ;
  assign wci_reqERR_5$EN =
	     WILL_FIRE_RL_wci_wrkBusy_5 &&
	     wci_wciResponse_5$wget[33:32] == 2'd3 &&
	     (wci_reqPend_5 == 2'd1 || wci_reqPend_5 == 2'd2 ||
	      wci_reqPend_5 == 2'd3) ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_F_T_T_T ;

  // register wci_reqERR_6
  assign wci_reqERR_6$D_IN =
	     MUX_wci_reqERR_6$write_1__SEL_1 ?
	       MUX_wci_reqERR_6$write_1__VAL_1 :
	       3'd0 ;
  assign wci_reqERR_6$EN =
	     WILL_FIRE_RL_wci_wrkBusy_6 &&
	     wci_wciResponse_6$wget[33:32] == 2'd3 &&
	     (wci_reqPend_6 == 2'd1 || wci_reqPend_6 == 2'd2 ||
	      wci_reqPend_6 == 2'd3) ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_F_T_T_T ;

  // register wci_reqERR_7
  assign wci_reqERR_7$D_IN =
	     MUX_wci_reqERR_7$write_1__SEL_1 ?
	       MUX_wci_reqERR_7$write_1__VAL_1 :
	       3'd0 ;
  assign wci_reqERR_7$EN =
	     WILL_FIRE_RL_wci_wrkBusy_7 &&
	     wci_wciResponse_7$wget[33:32] == 2'd3 &&
	     (wci_reqPend_7 == 2'd1 || wci_reqPend_7 == 2'd2 ||
	      wci_reqPend_7 == 2'd3) ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_F_T_T_T ;

  // register wci_reqERR_8
  assign wci_reqERR_8$D_IN =
	     MUX_wci_reqERR_8$write_1__SEL_1 ?
	       MUX_wci_reqERR_8$write_1__VAL_1 :
	       3'd0 ;
  assign wci_reqERR_8$EN =
	     WILL_FIRE_RL_wci_wrkBusy_8 &&
	     wci_wciResponse_8$wget[33:32] == 2'd3 &&
	     (wci_reqPend_8 == 2'd1 || wci_reqPend_8 == 2'd2 ||
	      wci_reqPend_8 == 2'd3) ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_F_T_T_T ;

  // register wci_reqERR_9
  assign wci_reqERR_9$D_IN =
	     MUX_wci_reqERR_9$write_1__SEL_1 ?
	       MUX_wci_reqERR_9$write_1__VAL_1 :
	       3'd0 ;
  assign wci_reqERR_9$EN =
	     WILL_FIRE_RL_wci_wrkBusy_9 &&
	     wci_wciResponse_9$wget[33:32] == 2'd3 &&
	     (wci_reqPend_9 == 2'd1 || wci_reqPend_9 == 2'd2 ||
	      wci_reqPend_9 == 2'd3) ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T ;

  // register wci_reqFAIL
  assign wci_reqFAIL$D_IN =
	     MUX_wci_reqFAIL$write_1__SEL_1 ?
	       MUX_wci_reqFAIL$write_1__VAL_1 :
	       3'd0 ;
  assign wci_reqFAIL$EN =
	     WILL_FIRE_RL_wci_wrkBusy &&
	     wci_wciResponse$wget[33:32] == 2'd2 &&
	     (wci_reqPend == 2'd1 || wci_reqPend == 2'd2 ||
	      wci_reqPend == 2'd3) ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_T_F_F_T_T_T ;

  // register wci_reqFAIL_1
  assign wci_reqFAIL_1$D_IN =
	     MUX_wci_reqFAIL_1$write_1__SEL_1 ?
	       MUX_wci_reqFAIL_1$write_1__VAL_1 :
	       3'd0 ;
  assign wci_reqFAIL_1$EN =
	     WILL_FIRE_RL_wci_wrkBusy_1 &&
	     wci_wciResponse_1$wget[33:32] == 2'd2 &&
	     (wci_reqPend_1 == 2'd1 || wci_reqPend_1 == 2'd2 ||
	      wci_reqPend_1 == 2'd3) ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_T_F_F_T_T_T ;

  // register wci_reqFAIL_10
  assign wci_reqFAIL_10$D_IN =
	     MUX_wci_reqFAIL_10$write_1__SEL_1 ?
	       MUX_wci_reqFAIL_10$write_1__VAL_1 :
	       3'd0 ;
  assign wci_reqFAIL_10$EN =
	     WILL_FIRE_RL_wci_wrkBusy_10 &&
	     wci_wciResponse_10$wget[33:32] == 2'd2 &&
	     (wci_reqPend_10 == 2'd1 || wci_reqPend_10 == 2'd2 ||
	      wci_reqPend_10 == 2'd3) ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T ;

  // register wci_reqFAIL_11
  assign wci_reqFAIL_11$D_IN =
	     MUX_wci_reqFAIL_11$write_1__SEL_1 ?
	       MUX_wci_reqFAIL_11$write_1__VAL_1 :
	       3'd0 ;
  assign wci_reqFAIL_11$EN =
	     WILL_FIRE_RL_wci_wrkBusy_11 &&
	     wci_wciResponse_11$wget[33:32] == 2'd2 &&
	     (wci_reqPend_11 == 2'd1 || wci_reqPend_11 == 2'd2 ||
	      wci_reqPend_11 == 2'd3) ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T ;

  // register wci_reqFAIL_12
  assign wci_reqFAIL_12$D_IN =
	     MUX_wci_reqFAIL_12$write_1__SEL_1 ?
	       MUX_wci_reqFAIL_12$write_1__VAL_1 :
	       3'd0 ;
  assign wci_reqFAIL_12$EN =
	     WILL_FIRE_RL_wci_wrkBusy_12 &&
	     wci_wciResponse_12$wget[33:32] == 2'd2 &&
	     (wci_reqPend_12 == 2'd1 || wci_reqPend_12 == 2'd2 ||
	      wci_reqPend_12 == 2'd3) ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T ;

  // register wci_reqFAIL_13
  assign wci_reqFAIL_13$D_IN =
	     MUX_wci_reqFAIL_13$write_1__SEL_1 ?
	       MUX_wci_reqFAIL_13$write_1__VAL_1 :
	       3'd0 ;
  assign wci_reqFAIL_13$EN =
	     WILL_FIRE_RL_wci_wrkBusy_13 &&
	     wci_wciResponse_13$wget[33:32] == 2'd2 &&
	     (wci_reqPend_13 == 2'd1 || wci_reqPend_13 == 2'd2 ||
	      wci_reqPend_13 == 2'd3) ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T ;

  // register wci_reqFAIL_14
  assign wci_reqFAIL_14$D_IN =
	     MUX_wci_reqFAIL_14$write_1__SEL_1 ?
	       MUX_wci_reqFAIL_14$write_1__VAL_1 :
	       3'd0 ;
  assign wci_reqFAIL_14$EN =
	     WILL_FIRE_RL_wci_wrkBusy_14 &&
	     wci_wciResponse_14$wget[33:32] == 2'd2 &&
	     (wci_reqPend_14 == 2'd1 || wci_reqPend_14 == 2'd2 ||
	      wci_reqPend_14 == 2'd3) ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T ;

  // register wci_reqFAIL_2
  assign wci_reqFAIL_2$D_IN =
	     MUX_wci_reqFAIL_2$write_1__SEL_1 ?
	       MUX_wci_reqFAIL_2$write_1__VAL_1 :
	       3'd0 ;
  assign wci_reqFAIL_2$EN =
	     WILL_FIRE_RL_wci_wrkBusy_2 &&
	     wci_wciResponse_2$wget[33:32] == 2'd2 &&
	     (wci_reqPend_2 == 2'd1 || wci_reqPend_2 == 2'd2 ||
	      wci_reqPend_2 == 2'd3) ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_F_F_T_T_T ;

  // register wci_reqFAIL_3
  assign wci_reqFAIL_3$D_IN =
	     MUX_wci_reqFAIL_3$write_1__SEL_1 ?
	       MUX_wci_reqFAIL_3$write_1__VAL_1 :
	       3'd0 ;
  assign wci_reqFAIL_3$EN =
	     WILL_FIRE_RL_wci_wrkBusy_3 &&
	     wci_wciResponse_3$wget[33:32] == 2'd2 &&
	     (wci_reqPend_3 == 2'd1 || wci_reqPend_3 == 2'd2 ||
	      wci_reqPend_3 == 2'd3) ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_F_F_T_T_T ;

  // register wci_reqFAIL_4
  assign wci_reqFAIL_4$D_IN =
	     MUX_wci_reqFAIL_4$write_1__SEL_1 ?
	       MUX_wci_reqFAIL_4$write_1__VAL_1 :
	       3'd0 ;
  assign wci_reqFAIL_4$EN =
	     WILL_FIRE_RL_wci_wrkBusy_4 &&
	     wci_wciResponse_4$wget[33:32] == 2'd2 &&
	     (wci_reqPend_4 == 2'd1 || wci_reqPend_4 == 2'd2 ||
	      wci_reqPend_4 == 2'd3) ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_F_F_T_T_T ;

  // register wci_reqFAIL_5
  assign wci_reqFAIL_5$D_IN =
	     MUX_wci_reqFAIL_5$write_1__SEL_1 ?
	       MUX_wci_reqFAIL_5$write_1__VAL_1 :
	       3'd0 ;
  assign wci_reqFAIL_5$EN =
	     WILL_FIRE_RL_wci_wrkBusy_5 &&
	     wci_wciResponse_5$wget[33:32] == 2'd2 &&
	     (wci_reqPend_5 == 2'd1 || wci_reqPend_5 == 2'd2 ||
	      wci_reqPend_5 == 2'd3) ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_F_T_T_T ;

  // register wci_reqFAIL_6
  assign wci_reqFAIL_6$D_IN =
	     MUX_wci_reqFAIL_6$write_1__SEL_1 ?
	       MUX_wci_reqFAIL_6$write_1__VAL_1 :
	       3'd0 ;
  assign wci_reqFAIL_6$EN =
	     WILL_FIRE_RL_wci_wrkBusy_6 &&
	     wci_wciResponse_6$wget[33:32] == 2'd2 &&
	     (wci_reqPend_6 == 2'd1 || wci_reqPend_6 == 2'd2 ||
	      wci_reqPend_6 == 2'd3) ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_F_T_T_T ;

  // register wci_reqFAIL_7
  assign wci_reqFAIL_7$D_IN =
	     MUX_wci_reqFAIL_7$write_1__SEL_1 ?
	       MUX_wci_reqFAIL_7$write_1__VAL_1 :
	       3'd0 ;
  assign wci_reqFAIL_7$EN =
	     WILL_FIRE_RL_wci_wrkBusy_7 &&
	     wci_wciResponse_7$wget[33:32] == 2'd2 &&
	     (wci_reqPend_7 == 2'd1 || wci_reqPend_7 == 2'd2 ||
	      wci_reqPend_7 == 2'd3) ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_F_T_T_T ;

  // register wci_reqFAIL_8
  assign wci_reqFAIL_8$D_IN =
	     MUX_wci_reqFAIL_8$write_1__SEL_1 ?
	       MUX_wci_reqFAIL_8$write_1__VAL_1 :
	       3'd0 ;
  assign wci_reqFAIL_8$EN =
	     WILL_FIRE_RL_wci_wrkBusy_8 &&
	     wci_wciResponse_8$wget[33:32] == 2'd2 &&
	     (wci_reqPend_8 == 2'd1 || wci_reqPend_8 == 2'd2 ||
	      wci_reqPend_8 == 2'd3) ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_F_T_T_T ;

  // register wci_reqFAIL_9
  assign wci_reqFAIL_9$D_IN =
	     MUX_wci_reqFAIL_9$write_1__SEL_1 ?
	       MUX_wci_reqFAIL_9$write_1__VAL_1 :
	       3'd0 ;
  assign wci_reqFAIL_9$EN =
	     WILL_FIRE_RL_wci_wrkBusy_9 &&
	     wci_wciResponse_9$wget[33:32] == 2'd2 &&
	     (wci_reqPend_9 == 2'd1 || wci_reqPend_9 == 2'd2 ||
	      wci_reqPend_9 == 2'd3) ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T ;

  // register wci_reqF_10_c_r
  assign wci_reqF_10_c_r$D_IN =
	     WILL_FIRE_RL_wci_reqF_10_incCtr ?
	       MUX_wci_reqF_10_c_r$write_1__VAL_1 :
	       MUX_wci_reqF_10_c_r$write_1__VAL_2 ;
  assign wci_reqF_10_c_r$EN =
	     WILL_FIRE_RL_wci_reqF_10_incCtr ||
	     WILL_FIRE_RL_wci_reqF_10_decCtr ;

  // register wci_reqF_10_q_0
  always@(MUX_wci_reqF_10_q_0$write_1__SEL_1 or
	  MUX_wci_reqF_10_q_0$write_1__VAL_1 or
	  WILL_FIRE_RL_wci_reqF_10_both or
	  MUX_wci_reqF_10_q_0$write_1__VAL_2 or
	  WILL_FIRE_RL_wci_reqF_10_decCtr)
  begin
    case (1'b1) // synopsys parallel_case
      MUX_wci_reqF_10_q_0$write_1__SEL_1:
	  wci_reqF_10_q_0$D_IN = MUX_wci_reqF_10_q_0$write_1__VAL_1;
      WILL_FIRE_RL_wci_reqF_10_both:
	  wci_reqF_10_q_0$D_IN = MUX_wci_reqF_10_q_0$write_1__VAL_2;
      WILL_FIRE_RL_wci_reqF_10_decCtr:
	  wci_reqF_10_q_0$D_IN = 72'h0000000000AAAAAAAA;
      default: wci_reqF_10_q_0$D_IN =
		   72'hAAAAAAAAAAAAAAAAAA /* unspecified value */ ;
    endcase
  end
  assign wci_reqF_10_q_0$EN =
	     WILL_FIRE_RL_wci_reqF_10_incCtr && !wci_reqF_10_c_r ||
	     WILL_FIRE_RL_wci_reqF_10_both ||
	     WILL_FIRE_RL_wci_reqF_10_decCtr ;

  // register wci_reqF_11_c_r
  assign wci_reqF_11_c_r$D_IN =
	     WILL_FIRE_RL_wci_reqF_11_incCtr ?
	       MUX_wci_reqF_11_c_r$write_1__VAL_1 :
	       MUX_wci_reqF_11_c_r$write_1__VAL_2 ;
  assign wci_reqF_11_c_r$EN =
	     WILL_FIRE_RL_wci_reqF_11_incCtr ||
	     WILL_FIRE_RL_wci_reqF_11_decCtr ;

  // register wci_reqF_11_q_0
  always@(MUX_wci_reqF_11_q_0$write_1__SEL_1 or
	  MUX_wci_reqF_11_q_0$write_1__VAL_1 or
	  WILL_FIRE_RL_wci_reqF_11_both or
	  MUX_wci_reqF_11_q_0$write_1__VAL_2 or
	  WILL_FIRE_RL_wci_reqF_11_decCtr)
  begin
    case (1'b1) // synopsys parallel_case
      MUX_wci_reqF_11_q_0$write_1__SEL_1:
	  wci_reqF_11_q_0$D_IN = MUX_wci_reqF_11_q_0$write_1__VAL_1;
      WILL_FIRE_RL_wci_reqF_11_both:
	  wci_reqF_11_q_0$D_IN = MUX_wci_reqF_11_q_0$write_1__VAL_2;
      WILL_FIRE_RL_wci_reqF_11_decCtr:
	  wci_reqF_11_q_0$D_IN = 72'h0000000000AAAAAAAA;
      default: wci_reqF_11_q_0$D_IN =
		   72'hAAAAAAAAAAAAAAAAAA /* unspecified value */ ;
    endcase
  end
  assign wci_reqF_11_q_0$EN =
	     WILL_FIRE_RL_wci_reqF_11_incCtr && !wci_reqF_11_c_r ||
	     WILL_FIRE_RL_wci_reqF_11_both ||
	     WILL_FIRE_RL_wci_reqF_11_decCtr ;

  // register wci_reqF_12_c_r
  assign wci_reqF_12_c_r$D_IN =
	     WILL_FIRE_RL_wci_reqF_12_incCtr ?
	       MUX_wci_reqF_12_c_r$write_1__VAL_1 :
	       MUX_wci_reqF_12_c_r$write_1__VAL_2 ;
  assign wci_reqF_12_c_r$EN =
	     WILL_FIRE_RL_wci_reqF_12_incCtr ||
	     WILL_FIRE_RL_wci_reqF_12_decCtr ;

  // register wci_reqF_12_q_0
  always@(MUX_wci_reqF_12_q_0$write_1__SEL_1 or
	  MUX_wci_reqF_12_q_0$write_1__VAL_1 or
	  WILL_FIRE_RL_wci_reqF_12_both or
	  MUX_wci_reqF_12_q_0$write_1__VAL_2 or
	  WILL_FIRE_RL_wci_reqF_12_decCtr)
  begin
    case (1'b1) // synopsys parallel_case
      MUX_wci_reqF_12_q_0$write_1__SEL_1:
	  wci_reqF_12_q_0$D_IN = MUX_wci_reqF_12_q_0$write_1__VAL_1;
      WILL_FIRE_RL_wci_reqF_12_both:
	  wci_reqF_12_q_0$D_IN = MUX_wci_reqF_12_q_0$write_1__VAL_2;
      WILL_FIRE_RL_wci_reqF_12_decCtr:
	  wci_reqF_12_q_0$D_IN = 72'h0000000000AAAAAAAA;
      default: wci_reqF_12_q_0$D_IN =
		   72'hAAAAAAAAAAAAAAAAAA /* unspecified value */ ;
    endcase
  end
  assign wci_reqF_12_q_0$EN =
	     WILL_FIRE_RL_wci_reqF_12_incCtr && !wci_reqF_12_c_r ||
	     WILL_FIRE_RL_wci_reqF_12_both ||
	     WILL_FIRE_RL_wci_reqF_12_decCtr ;

  // register wci_reqF_13_c_r
  assign wci_reqF_13_c_r$D_IN =
	     WILL_FIRE_RL_wci_reqF_13_incCtr ?
	       MUX_wci_reqF_13_c_r$write_1__VAL_1 :
	       MUX_wci_reqF_13_c_r$write_1__VAL_2 ;
  assign wci_reqF_13_c_r$EN =
	     WILL_FIRE_RL_wci_reqF_13_incCtr ||
	     WILL_FIRE_RL_wci_reqF_13_decCtr ;

  // register wci_reqF_13_q_0
  always@(MUX_wci_reqF_13_q_0$write_1__SEL_1 or
	  MUX_wci_reqF_13_q_0$write_1__VAL_1 or
	  WILL_FIRE_RL_wci_reqF_13_both or
	  MUX_wci_reqF_13_q_0$write_1__VAL_2 or
	  WILL_FIRE_RL_wci_reqF_13_decCtr)
  begin
    case (1'b1) // synopsys parallel_case
      MUX_wci_reqF_13_q_0$write_1__SEL_1:
	  wci_reqF_13_q_0$D_IN = MUX_wci_reqF_13_q_0$write_1__VAL_1;
      WILL_FIRE_RL_wci_reqF_13_both:
	  wci_reqF_13_q_0$D_IN = MUX_wci_reqF_13_q_0$write_1__VAL_2;
      WILL_FIRE_RL_wci_reqF_13_decCtr:
	  wci_reqF_13_q_0$D_IN = 72'h0000000000AAAAAAAA;
      default: wci_reqF_13_q_0$D_IN =
		   72'hAAAAAAAAAAAAAAAAAA /* unspecified value */ ;
    endcase
  end
  assign wci_reqF_13_q_0$EN =
	     WILL_FIRE_RL_wci_reqF_13_incCtr && !wci_reqF_13_c_r ||
	     WILL_FIRE_RL_wci_reqF_13_both ||
	     WILL_FIRE_RL_wci_reqF_13_decCtr ;

  // register wci_reqF_14_c_r
  assign wci_reqF_14_c_r$D_IN =
	     WILL_FIRE_RL_wci_reqF_14_incCtr ?
	       MUX_wci_reqF_14_c_r$write_1__VAL_1 :
	       MUX_wci_reqF_14_c_r$write_1__VAL_2 ;
  assign wci_reqF_14_c_r$EN =
	     WILL_FIRE_RL_wci_reqF_14_incCtr ||
	     WILL_FIRE_RL_wci_reqF_14_decCtr ;

  // register wci_reqF_14_q_0
  always@(MUX_wci_reqF_14_q_0$write_1__SEL_1 or
	  MUX_wci_reqF_14_q_0$write_1__VAL_1 or
	  WILL_FIRE_RL_wci_reqF_14_both or
	  MUX_wci_reqF_14_q_0$write_1__VAL_2 or
	  WILL_FIRE_RL_wci_reqF_14_decCtr)
  begin
    case (1'b1) // synopsys parallel_case
      MUX_wci_reqF_14_q_0$write_1__SEL_1:
	  wci_reqF_14_q_0$D_IN = MUX_wci_reqF_14_q_0$write_1__VAL_1;
      WILL_FIRE_RL_wci_reqF_14_both:
	  wci_reqF_14_q_0$D_IN = MUX_wci_reqF_14_q_0$write_1__VAL_2;
      WILL_FIRE_RL_wci_reqF_14_decCtr:
	  wci_reqF_14_q_0$D_IN = 72'h0000000000AAAAAAAA;
      default: wci_reqF_14_q_0$D_IN =
		   72'hAAAAAAAAAAAAAAAAAA /* unspecified value */ ;
    endcase
  end
  assign wci_reqF_14_q_0$EN =
	     WILL_FIRE_RL_wci_reqF_14_incCtr && !wci_reqF_14_c_r ||
	     WILL_FIRE_RL_wci_reqF_14_both ||
	     WILL_FIRE_RL_wci_reqF_14_decCtr ;

  // register wci_reqF_1_c_r
  assign wci_reqF_1_c_r$D_IN =
	     WILL_FIRE_RL_wci_reqF_1_incCtr ?
	       MUX_wci_reqF_1_c_r$write_1__VAL_1 :
	       MUX_wci_reqF_1_c_r$write_1__VAL_2 ;
  assign wci_reqF_1_c_r$EN =
	     WILL_FIRE_RL_wci_reqF_1_incCtr ||
	     WILL_FIRE_RL_wci_reqF_1_decCtr ;

  // register wci_reqF_1_q_0
  always@(WILL_FIRE_RL_wci_reqF_1_both or
	  MUX_wci_reqF_1_q_0$write_1__VAL_1 or
	  MUX_wci_reqF_1_q_0$write_1__SEL_2 or
	  MUX_wci_reqF_1_q_0$write_1__VAL_2 or WILL_FIRE_RL_wci_reqF_1_decCtr)
  begin
    case (1'b1) // synopsys parallel_case
      WILL_FIRE_RL_wci_reqF_1_both:
	  wci_reqF_1_q_0$D_IN = MUX_wci_reqF_1_q_0$write_1__VAL_1;
      MUX_wci_reqF_1_q_0$write_1__SEL_2:
	  wci_reqF_1_q_0$D_IN = MUX_wci_reqF_1_q_0$write_1__VAL_2;
      WILL_FIRE_RL_wci_reqF_1_decCtr:
	  wci_reqF_1_q_0$D_IN = 72'h0000000000AAAAAAAA;
      default: wci_reqF_1_q_0$D_IN =
		   72'hAAAAAAAAAAAAAAAAAA /* unspecified value */ ;
    endcase
  end
  assign wci_reqF_1_q_0$EN =
	     WILL_FIRE_RL_wci_reqF_1_both ||
	     WILL_FIRE_RL_wci_reqF_1_incCtr && !wci_reqF_1_c_r ||
	     WILL_FIRE_RL_wci_reqF_1_decCtr ;

  // register wci_reqF_2_c_r
  assign wci_reqF_2_c_r$D_IN =
	     WILL_FIRE_RL_wci_reqF_2_incCtr ?
	       MUX_wci_reqF_2_c_r$write_1__VAL_1 :
	       MUX_wci_reqF_2_c_r$write_1__VAL_2 ;
  assign wci_reqF_2_c_r$EN =
	     WILL_FIRE_RL_wci_reqF_2_incCtr ||
	     WILL_FIRE_RL_wci_reqF_2_decCtr ;

  // register wci_reqF_2_q_0
  always@(WILL_FIRE_RL_wci_reqF_2_both or
	  MUX_wci_reqF_2_q_0$write_1__VAL_1 or
	  MUX_wci_reqF_2_q_0$write_1__SEL_2 or
	  MUX_wci_reqF_2_q_0$write_1__VAL_2 or WILL_FIRE_RL_wci_reqF_2_decCtr)
  begin
    case (1'b1) // synopsys parallel_case
      WILL_FIRE_RL_wci_reqF_2_both:
	  wci_reqF_2_q_0$D_IN = MUX_wci_reqF_2_q_0$write_1__VAL_1;
      MUX_wci_reqF_2_q_0$write_1__SEL_2:
	  wci_reqF_2_q_0$D_IN = MUX_wci_reqF_2_q_0$write_1__VAL_2;
      WILL_FIRE_RL_wci_reqF_2_decCtr:
	  wci_reqF_2_q_0$D_IN = 72'h0000000000AAAAAAAA;
      default: wci_reqF_2_q_0$D_IN =
		   72'hAAAAAAAAAAAAAAAAAA /* unspecified value */ ;
    endcase
  end
  assign wci_reqF_2_q_0$EN =
	     WILL_FIRE_RL_wci_reqF_2_both ||
	     WILL_FIRE_RL_wci_reqF_2_incCtr && !wci_reqF_2_c_r ||
	     WILL_FIRE_RL_wci_reqF_2_decCtr ;

  // register wci_reqF_3_c_r
  assign wci_reqF_3_c_r$D_IN =
	     WILL_FIRE_RL_wci_reqF_3_incCtr ?
	       MUX_wci_reqF_3_c_r$write_1__VAL_1 :
	       MUX_wci_reqF_3_c_r$write_1__VAL_2 ;
  assign wci_reqF_3_c_r$EN =
	     WILL_FIRE_RL_wci_reqF_3_incCtr ||
	     WILL_FIRE_RL_wci_reqF_3_decCtr ;

  // register wci_reqF_3_q_0
  always@(WILL_FIRE_RL_wci_reqF_3_both or
	  MUX_wci_reqF_3_q_0$write_1__VAL_1 or
	  MUX_wci_reqF_3_q_0$write_1__SEL_2 or
	  MUX_wci_reqF_3_q_0$write_1__VAL_2 or WILL_FIRE_RL_wci_reqF_3_decCtr)
  begin
    case (1'b1) // synopsys parallel_case
      WILL_FIRE_RL_wci_reqF_3_both:
	  wci_reqF_3_q_0$D_IN = MUX_wci_reqF_3_q_0$write_1__VAL_1;
      MUX_wci_reqF_3_q_0$write_1__SEL_2:
	  wci_reqF_3_q_0$D_IN = MUX_wci_reqF_3_q_0$write_1__VAL_2;
      WILL_FIRE_RL_wci_reqF_3_decCtr:
	  wci_reqF_3_q_0$D_IN = 72'h0000000000AAAAAAAA;
      default: wci_reqF_3_q_0$D_IN =
		   72'hAAAAAAAAAAAAAAAAAA /* unspecified value */ ;
    endcase
  end
  assign wci_reqF_3_q_0$EN =
	     WILL_FIRE_RL_wci_reqF_3_both ||
	     WILL_FIRE_RL_wci_reqF_3_incCtr && !wci_reqF_3_c_r ||
	     WILL_FIRE_RL_wci_reqF_3_decCtr ;

  // register wci_reqF_4_c_r
  assign wci_reqF_4_c_r$D_IN =
	     WILL_FIRE_RL_wci_reqF_4_incCtr ?
	       MUX_wci_reqF_4_c_r$write_1__VAL_1 :
	       MUX_wci_reqF_4_c_r$write_1__VAL_2 ;
  assign wci_reqF_4_c_r$EN =
	     WILL_FIRE_RL_wci_reqF_4_incCtr ||
	     WILL_FIRE_RL_wci_reqF_4_decCtr ;

  // register wci_reqF_4_q_0
  always@(WILL_FIRE_RL_wci_reqF_4_both or
	  MUX_wci_reqF_4_q_0$write_1__VAL_1 or
	  MUX_wci_reqF_4_q_0$write_1__SEL_2 or
	  MUX_wci_reqF_4_q_0$write_1__VAL_2 or WILL_FIRE_RL_wci_reqF_4_decCtr)
  begin
    case (1'b1) // synopsys parallel_case
      WILL_FIRE_RL_wci_reqF_4_both:
	  wci_reqF_4_q_0$D_IN = MUX_wci_reqF_4_q_0$write_1__VAL_1;
      MUX_wci_reqF_4_q_0$write_1__SEL_2:
	  wci_reqF_4_q_0$D_IN = MUX_wci_reqF_4_q_0$write_1__VAL_2;
      WILL_FIRE_RL_wci_reqF_4_decCtr:
	  wci_reqF_4_q_0$D_IN = 72'h0000000000AAAAAAAA;
      default: wci_reqF_4_q_0$D_IN =
		   72'hAAAAAAAAAAAAAAAAAA /* unspecified value */ ;
    endcase
  end
  assign wci_reqF_4_q_0$EN =
	     WILL_FIRE_RL_wci_reqF_4_both ||
	     WILL_FIRE_RL_wci_reqF_4_incCtr && !wci_reqF_4_c_r ||
	     WILL_FIRE_RL_wci_reqF_4_decCtr ;

  // register wci_reqF_5_c_r
  assign wci_reqF_5_c_r$D_IN =
	     WILL_FIRE_RL_wci_reqF_5_incCtr ?
	       MUX_wci_reqF_5_c_r$write_1__VAL_1 :
	       MUX_wci_reqF_5_c_r$write_1__VAL_2 ;
  assign wci_reqF_5_c_r$EN =
	     WILL_FIRE_RL_wci_reqF_5_incCtr ||
	     WILL_FIRE_RL_wci_reqF_5_decCtr ;

  // register wci_reqF_5_q_0
  always@(WILL_FIRE_RL_wci_reqF_5_both or
	  MUX_wci_reqF_5_q_0$write_1__VAL_1 or
	  MUX_wci_reqF_5_q_0$write_1__SEL_2 or
	  MUX_wci_reqF_5_q_0$write_1__VAL_2 or WILL_FIRE_RL_wci_reqF_5_decCtr)
  begin
    case (1'b1) // synopsys parallel_case
      WILL_FIRE_RL_wci_reqF_5_both:
	  wci_reqF_5_q_0$D_IN = MUX_wci_reqF_5_q_0$write_1__VAL_1;
      MUX_wci_reqF_5_q_0$write_1__SEL_2:
	  wci_reqF_5_q_0$D_IN = MUX_wci_reqF_5_q_0$write_1__VAL_2;
      WILL_FIRE_RL_wci_reqF_5_decCtr:
	  wci_reqF_5_q_0$D_IN = 72'h0000000000AAAAAAAA;
      default: wci_reqF_5_q_0$D_IN =
		   72'hAAAAAAAAAAAAAAAAAA /* unspecified value */ ;
    endcase
  end
  assign wci_reqF_5_q_0$EN =
	     WILL_FIRE_RL_wci_reqF_5_both ||
	     WILL_FIRE_RL_wci_reqF_5_incCtr && !wci_reqF_5_c_r ||
	     WILL_FIRE_RL_wci_reqF_5_decCtr ;

  // register wci_reqF_6_c_r
  assign wci_reqF_6_c_r$D_IN =
	     WILL_FIRE_RL_wci_reqF_6_incCtr ?
	       MUX_wci_reqF_6_c_r$write_1__VAL_1 :
	       MUX_wci_reqF_6_c_r$write_1__VAL_2 ;
  assign wci_reqF_6_c_r$EN =
	     WILL_FIRE_RL_wci_reqF_6_incCtr ||
	     WILL_FIRE_RL_wci_reqF_6_decCtr ;

  // register wci_reqF_6_q_0
  always@(WILL_FIRE_RL_wci_reqF_6_both or
	  MUX_wci_reqF_6_q_0$write_1__VAL_1 or
	  MUX_wci_reqF_6_q_0$write_1__SEL_2 or
	  MUX_wci_reqF_6_q_0$write_1__VAL_2 or WILL_FIRE_RL_wci_reqF_6_decCtr)
  begin
    case (1'b1) // synopsys parallel_case
      WILL_FIRE_RL_wci_reqF_6_both:
	  wci_reqF_6_q_0$D_IN = MUX_wci_reqF_6_q_0$write_1__VAL_1;
      MUX_wci_reqF_6_q_0$write_1__SEL_2:
	  wci_reqF_6_q_0$D_IN = MUX_wci_reqF_6_q_0$write_1__VAL_2;
      WILL_FIRE_RL_wci_reqF_6_decCtr:
	  wci_reqF_6_q_0$D_IN = 72'h0000000000AAAAAAAA;
      default: wci_reqF_6_q_0$D_IN =
		   72'hAAAAAAAAAAAAAAAAAA /* unspecified value */ ;
    endcase
  end
  assign wci_reqF_6_q_0$EN =
	     WILL_FIRE_RL_wci_reqF_6_both ||
	     WILL_FIRE_RL_wci_reqF_6_incCtr && !wci_reqF_6_c_r ||
	     WILL_FIRE_RL_wci_reqF_6_decCtr ;

  // register wci_reqF_7_c_r
  assign wci_reqF_7_c_r$D_IN =
	     WILL_FIRE_RL_wci_reqF_7_incCtr ?
	       MUX_wci_reqF_7_c_r$write_1__VAL_1 :
	       MUX_wci_reqF_7_c_r$write_1__VAL_2 ;
  assign wci_reqF_7_c_r$EN =
	     WILL_FIRE_RL_wci_reqF_7_incCtr ||
	     WILL_FIRE_RL_wci_reqF_7_decCtr ;

  // register wci_reqF_7_q_0
  always@(WILL_FIRE_RL_wci_reqF_7_both or
	  MUX_wci_reqF_7_q_0$write_1__VAL_1 or
	  MUX_wci_reqF_7_q_0$write_1__SEL_2 or
	  MUX_wci_reqF_7_q_0$write_1__VAL_2 or WILL_FIRE_RL_wci_reqF_7_decCtr)
  begin
    case (1'b1) // synopsys parallel_case
      WILL_FIRE_RL_wci_reqF_7_both:
	  wci_reqF_7_q_0$D_IN = MUX_wci_reqF_7_q_0$write_1__VAL_1;
      MUX_wci_reqF_7_q_0$write_1__SEL_2:
	  wci_reqF_7_q_0$D_IN = MUX_wci_reqF_7_q_0$write_1__VAL_2;
      WILL_FIRE_RL_wci_reqF_7_decCtr:
	  wci_reqF_7_q_0$D_IN = 72'h0000000000AAAAAAAA;
      default: wci_reqF_7_q_0$D_IN =
		   72'hAAAAAAAAAAAAAAAAAA /* unspecified value */ ;
    endcase
  end
  assign wci_reqF_7_q_0$EN =
	     WILL_FIRE_RL_wci_reqF_7_both ||
	     WILL_FIRE_RL_wci_reqF_7_incCtr && !wci_reqF_7_c_r ||
	     WILL_FIRE_RL_wci_reqF_7_decCtr ;

  // register wci_reqF_8_c_r
  assign wci_reqF_8_c_r$D_IN =
	     WILL_FIRE_RL_wci_reqF_8_incCtr ?
	       MUX_wci_reqF_8_c_r$write_1__VAL_1 :
	       MUX_wci_reqF_8_c_r$write_1__VAL_2 ;
  assign wci_reqF_8_c_r$EN =
	     WILL_FIRE_RL_wci_reqF_8_incCtr ||
	     WILL_FIRE_RL_wci_reqF_8_decCtr ;

  // register wci_reqF_8_q_0
  always@(WILL_FIRE_RL_wci_reqF_8_both or
	  MUX_wci_reqF_8_q_0$write_1__VAL_1 or
	  MUX_wci_reqF_8_q_0$write_1__SEL_2 or
	  MUX_wci_reqF_8_q_0$write_1__VAL_2 or WILL_FIRE_RL_wci_reqF_8_decCtr)
  begin
    case (1'b1) // synopsys parallel_case
      WILL_FIRE_RL_wci_reqF_8_both:
	  wci_reqF_8_q_0$D_IN = MUX_wci_reqF_8_q_0$write_1__VAL_1;
      MUX_wci_reqF_8_q_0$write_1__SEL_2:
	  wci_reqF_8_q_0$D_IN = MUX_wci_reqF_8_q_0$write_1__VAL_2;
      WILL_FIRE_RL_wci_reqF_8_decCtr:
	  wci_reqF_8_q_0$D_IN = 72'h0000000000AAAAAAAA;
      default: wci_reqF_8_q_0$D_IN =
		   72'hAAAAAAAAAAAAAAAAAA /* unspecified value */ ;
    endcase
  end
  assign wci_reqF_8_q_0$EN =
	     WILL_FIRE_RL_wci_reqF_8_both ||
	     WILL_FIRE_RL_wci_reqF_8_incCtr && !wci_reqF_8_c_r ||
	     WILL_FIRE_RL_wci_reqF_8_decCtr ;

  // register wci_reqF_9_c_r
  assign wci_reqF_9_c_r$D_IN =
	     WILL_FIRE_RL_wci_reqF_9_incCtr ?
	       MUX_wci_reqF_9_c_r$write_1__VAL_1 :
	       MUX_wci_reqF_9_c_r$write_1__VAL_2 ;
  assign wci_reqF_9_c_r$EN =
	     WILL_FIRE_RL_wci_reqF_9_incCtr ||
	     WILL_FIRE_RL_wci_reqF_9_decCtr ;

  // register wci_reqF_9_q_0
  always@(WILL_FIRE_RL_wci_reqF_9_both or
	  MUX_wci_reqF_9_q_0$write_1__VAL_1 or
	  MUX_wci_reqF_9_q_0$write_1__SEL_2 or
	  MUX_wci_reqF_9_q_0$write_1__VAL_2 or WILL_FIRE_RL_wci_reqF_9_decCtr)
  begin
    case (1'b1) // synopsys parallel_case
      WILL_FIRE_RL_wci_reqF_9_both:
	  wci_reqF_9_q_0$D_IN = MUX_wci_reqF_9_q_0$write_1__VAL_1;
      MUX_wci_reqF_9_q_0$write_1__SEL_2:
	  wci_reqF_9_q_0$D_IN = MUX_wci_reqF_9_q_0$write_1__VAL_2;
      WILL_FIRE_RL_wci_reqF_9_decCtr:
	  wci_reqF_9_q_0$D_IN = 72'h0000000000AAAAAAAA;
      default: wci_reqF_9_q_0$D_IN =
		   72'hAAAAAAAAAAAAAAAAAA /* unspecified value */ ;
    endcase
  end
  assign wci_reqF_9_q_0$EN =
	     WILL_FIRE_RL_wci_reqF_9_both ||
	     WILL_FIRE_RL_wci_reqF_9_incCtr && !wci_reqF_9_c_r ||
	     WILL_FIRE_RL_wci_reqF_9_decCtr ;

  // register wci_reqF_c_r
  assign wci_reqF_c_r$D_IN =
	     WILL_FIRE_RL_wci_reqF_incCtr ?
	       MUX_wci_reqF_c_r$write_1__VAL_1 :
	       MUX_wci_reqF_c_r$write_1__VAL_2 ;
  assign wci_reqF_c_r$EN =
	     WILL_FIRE_RL_wci_reqF_incCtr || WILL_FIRE_RL_wci_reqF_decCtr ;

  // register wci_reqF_q_0
  always@(WILL_FIRE_RL_wci_reqF_both or
	  MUX_wci_reqF_q_0$write_1__VAL_1 or
	  MUX_wci_reqF_q_0$write_1__SEL_2 or
	  MUX_wci_reqF_q_0$write_1__VAL_2 or WILL_FIRE_RL_wci_reqF_decCtr)
  begin
    case (1'b1) // synopsys parallel_case
      WILL_FIRE_RL_wci_reqF_both:
	  wci_reqF_q_0$D_IN = MUX_wci_reqF_q_0$write_1__VAL_1;
      MUX_wci_reqF_q_0$write_1__SEL_2:
	  wci_reqF_q_0$D_IN = MUX_wci_reqF_q_0$write_1__VAL_2;
      WILL_FIRE_RL_wci_reqF_decCtr:
	  wci_reqF_q_0$D_IN = 72'h0000000000AAAAAAAA;
      default: wci_reqF_q_0$D_IN =
		   72'hAAAAAAAAAAAAAAAAAA /* unspecified value */ ;
    endcase
  end
  assign wci_reqF_q_0$EN =
	     WILL_FIRE_RL_wci_reqF_both ||
	     WILL_FIRE_RL_wci_reqF_incCtr && !wci_reqF_c_r ||
	     WILL_FIRE_RL_wci_reqF_decCtr ;

  // register wci_reqPend
  always@(MUX_wci_reqPend$write_1__SEL_1 or
	  WILL_FIRE_RL_cpDispatch_F_F_T_T_T_T or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_T_T_T or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_T_F_T_T)
  begin
    case (1'b1) // synopsys parallel_case
      MUX_wci_reqPend$write_1__SEL_1: wci_reqPend$D_IN = 2'd0;
      WILL_FIRE_RL_cpDispatch_F_F_T_T_T_T: wci_reqPend$D_IN = 2'd1;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_T_T_T: wci_reqPend$D_IN = 2'd2;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_T_F_T_T: wci_reqPend$D_IN = 2'd3;
      default: wci_reqPend$D_IN = 2'b10 /* unspecified value */ ;
    endcase
  end
  assign wci_reqPend$EN =
	     WILL_FIRE_RL_wci_wrkBusy &&
	     wci_wciResponse$wget[33:32] != 2'd0 ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_T_F_T_T ;

  // register wci_reqPend_1
  always@(MUX_wci_reqPend_1$write_1__SEL_1 or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_T_T_T or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_T_T or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_F_T_T)
  begin
    case (1'b1) // synopsys parallel_case
      MUX_wci_reqPend_1$write_1__SEL_1: wci_reqPend_1$D_IN = 2'd0;
      WILL_FIRE_RL_cpDispatch_F_F_T_F_T_T_T: wci_reqPend_1$D_IN = 2'd1;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_T_T: wci_reqPend_1$D_IN = 2'd2;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_F_T_T: wci_reqPend_1$D_IN = 2'd3;
      default: wci_reqPend_1$D_IN = 2'b10 /* unspecified value */ ;
    endcase
  end
  assign wci_reqPend_1$EN =
	     WILL_FIRE_RL_wci_wrkBusy_1 &&
	     wci_wciResponse_1$wget[33:32] != 2'd0 ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_F_T_T ;

  // register wci_reqPend_10
  always@(MUX_wci_reqPend_10$write_1__SEL_1 or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_T_T or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T)
  begin
    case (1'b1) // synopsys parallel_case
      MUX_wci_reqPend_10$write_1__SEL_1: wci_reqPend_10$D_IN = 2'd0;
      WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_T_T:
	  wci_reqPend_10$D_IN = 2'd1;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T:
	  wci_reqPend_10$D_IN = 2'd2;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T:
	  wci_reqPend_10$D_IN = 2'd3;
      default: wci_reqPend_10$D_IN = 2'b10 /* unspecified value */ ;
    endcase
  end
  assign wci_reqPend_10$EN =
	     WILL_FIRE_RL_wci_wrkBusy_10 &&
	     wci_wciResponse_10$wget[33:32] != 2'd0 ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T ;

  // register wci_reqPend_11
  always@(MUX_wci_reqPend_11$write_1__SEL_1 or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_T_T or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T)
  begin
    case (1'b1) // synopsys parallel_case
      MUX_wci_reqPend_11$write_1__SEL_1: wci_reqPend_11$D_IN = 2'd0;
      WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_T_T:
	  wci_reqPend_11$D_IN = 2'd1;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T:
	  wci_reqPend_11$D_IN = 2'd2;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T:
	  wci_reqPend_11$D_IN = 2'd3;
      default: wci_reqPend_11$D_IN = 2'b10 /* unspecified value */ ;
    endcase
  end
  assign wci_reqPend_11$EN =
	     WILL_FIRE_RL_wci_wrkBusy_11 &&
	     wci_wciResponse_11$wget[33:32] != 2'd0 ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T ;

  // register wci_reqPend_12
  always@(MUX_wci_reqPend_12$write_1__SEL_1 or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T)
  begin
    case (1'b1) // synopsys parallel_case
      MUX_wci_reqPend_12$write_1__SEL_1: wci_reqPend_12$D_IN = 2'd0;
      WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T:
	  wci_reqPend_12$D_IN = 2'd1;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T:
	  wci_reqPend_12$D_IN = 2'd2;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T:
	  wci_reqPend_12$D_IN = 2'd3;
      default: wci_reqPend_12$D_IN = 2'b10 /* unspecified value */ ;
    endcase
  end
  assign wci_reqPend_12$EN =
	     WILL_FIRE_RL_wci_wrkBusy_12 &&
	     wci_wciResponse_12$wget[33:32] != 2'd0 ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T ;

  // register wci_reqPend_13
  always@(MUX_wci_reqPend_13$write_1__SEL_1 or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T)
  begin
    case (1'b1) // synopsys parallel_case
      MUX_wci_reqPend_13$write_1__SEL_1: wci_reqPend_13$D_IN = 2'd0;
      WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T:
	  wci_reqPend_13$D_IN = 2'd1;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T:
	  wci_reqPend_13$D_IN = 2'd2;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T:
	  wci_reqPend_13$D_IN = 2'd3;
      default: wci_reqPend_13$D_IN = 2'b10 /* unspecified value */ ;
    endcase
  end
  assign wci_reqPend_13$EN =
	     WILL_FIRE_RL_wci_wrkBusy_13 &&
	     wci_wciResponse_13$wget[33:32] != 2'd0 ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T ;

  // register wci_reqPend_14
  always@(MUX_wci_reqPend_14$write_1__SEL_1 or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T)
  begin
    case (1'b1) // synopsys parallel_case
      MUX_wci_reqPend_14$write_1__SEL_1: wci_reqPend_14$D_IN = 2'd0;
      WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T:
	  wci_reqPend_14$D_IN = 2'd1;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T:
	  wci_reqPend_14$D_IN = 2'd2;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T:
	  wci_reqPend_14$D_IN = 2'd3;
      default: wci_reqPend_14$D_IN = 2'b10 /* unspecified value */ ;
    endcase
  end
  assign wci_reqPend_14$EN =
	     WILL_FIRE_RL_wci_wrkBusy_14 &&
	     wci_wciResponse_14$wget[33:32] != 2'd0 ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T ;

  // register wci_reqPend_2
  always@(MUX_wci_reqPend_2$write_1__SEL_1 or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_T_T or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_T_T or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_F_T_T)
  begin
    case (1'b1) // synopsys parallel_case
      MUX_wci_reqPend_2$write_1__SEL_1: wci_reqPend_2$D_IN = 2'd0;
      WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_T_T: wci_reqPend_2$D_IN = 2'd1;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_T_T: wci_reqPend_2$D_IN = 2'd2;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_F_T_T: wci_reqPend_2$D_IN = 2'd3;
      default: wci_reqPend_2$D_IN = 2'b10 /* unspecified value */ ;
    endcase
  end
  assign wci_reqPend_2$EN =
	     WILL_FIRE_RL_wci_wrkBusy_2 &&
	     wci_wciResponse_2$wget[33:32] != 2'd0 ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_F_T_T ;

  // register wci_reqPend_3
  always@(MUX_wci_reqPend_3$write_1__SEL_1 or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_T_T or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_T_T or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_F_T_T)
  begin
    case (1'b1) // synopsys parallel_case
      MUX_wci_reqPend_3$write_1__SEL_1: wci_reqPend_3$D_IN = 2'd0;
      WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_T_T: wci_reqPend_3$D_IN = 2'd1;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_T_T: wci_reqPend_3$D_IN = 2'd2;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_F_T_T:
	  wci_reqPend_3$D_IN = 2'd3;
      default: wci_reqPend_3$D_IN = 2'b10 /* unspecified value */ ;
    endcase
  end
  assign wci_reqPend_3$EN =
	     WILL_FIRE_RL_wci_wrkBusy_3 &&
	     wci_wciResponse_3$wget[33:32] != 2'd0 ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_F_T_T ;

  // register wci_reqPend_4
  always@(MUX_wci_reqPend_4$write_1__SEL_1 or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_T_T or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_T_T or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_F_T_T)
  begin
    case (1'b1) // synopsys parallel_case
      MUX_wci_reqPend_4$write_1__SEL_1: wci_reqPend_4$D_IN = 2'd0;
      WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_T_T: wci_reqPend_4$D_IN = 2'd1;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_T_T:
	  wci_reqPend_4$D_IN = 2'd2;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_F_T_T:
	  wci_reqPend_4$D_IN = 2'd3;
      default: wci_reqPend_4$D_IN = 2'b10 /* unspecified value */ ;
    endcase
  end
  assign wci_reqPend_4$EN =
	     WILL_FIRE_RL_wci_wrkBusy_4 &&
	     wci_wciResponse_4$wget[33:32] != 2'd0 ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_F_T_T ;

  // register wci_reqPend_5
  always@(MUX_wci_reqPend_5$write_1__SEL_1 or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_T_T or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_T_T or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_F_T_T)
  begin
    case (1'b1) // synopsys parallel_case
      MUX_wci_reqPend_5$write_1__SEL_1: wci_reqPend_5$D_IN = 2'd0;
      WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_T_T:
	  wci_reqPend_5$D_IN = 2'd1;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_T_T:
	  wci_reqPend_5$D_IN = 2'd2;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_F_T_T:
	  wci_reqPend_5$D_IN = 2'd3;
      default: wci_reqPend_5$D_IN = 2'b10 /* unspecified value */ ;
    endcase
  end
  assign wci_reqPend_5$EN =
	     WILL_FIRE_RL_wci_wrkBusy_5 &&
	     wci_wciResponse_5$wget[33:32] != 2'd0 ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_F_T_T ;

  // register wci_reqPend_6
  always@(MUX_wci_reqPend_6$write_1__SEL_1 or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_T_T or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_T_T or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_F_T_T)
  begin
    case (1'b1) // synopsys parallel_case
      MUX_wci_reqPend_6$write_1__SEL_1: wci_reqPend_6$D_IN = 2'd0;
      WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_T_T:
	  wci_reqPend_6$D_IN = 2'd1;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_T_T:
	  wci_reqPend_6$D_IN = 2'd2;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_F_T_T:
	  wci_reqPend_6$D_IN = 2'd3;
      default: wci_reqPend_6$D_IN = 2'b10 /* unspecified value */ ;
    endcase
  end
  assign wci_reqPend_6$EN =
	     WILL_FIRE_RL_wci_wrkBusy_6 &&
	     wci_wciResponse_6$wget[33:32] != 2'd0 ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_F_T_T ;

  // register wci_reqPend_7
  always@(MUX_wci_reqPend_7$write_1__SEL_1 or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_T_T or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_T_T or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T)
  begin
    case (1'b1) // synopsys parallel_case
      MUX_wci_reqPend_7$write_1__SEL_1: wci_reqPend_7$D_IN = 2'd0;
      WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_T_T:
	  wci_reqPend_7$D_IN = 2'd1;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_T_T:
	  wci_reqPend_7$D_IN = 2'd2;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T:
	  wci_reqPend_7$D_IN = 2'd3;
      default: wci_reqPend_7$D_IN = 2'b10 /* unspecified value */ ;
    endcase
  end
  assign wci_reqPend_7$EN =
	     WILL_FIRE_RL_wci_wrkBusy_7 &&
	     wci_wciResponse_7$wget[33:32] != 2'd0 ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T ;

  // register wci_reqPend_8
  always@(MUX_wci_reqPend_8$write_1__SEL_1 or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_T_T or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T)
  begin
    case (1'b1) // synopsys parallel_case
      MUX_wci_reqPend_8$write_1__SEL_1: wci_reqPend_8$D_IN = 2'd0;
      WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_T_T:
	  wci_reqPend_8$D_IN = 2'd1;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T:
	  wci_reqPend_8$D_IN = 2'd2;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T:
	  wci_reqPend_8$D_IN = 2'd3;
      default: wci_reqPend_8$D_IN = 2'b10 /* unspecified value */ ;
    endcase
  end
  assign wci_reqPend_8$EN =
	     WILL_FIRE_RL_wci_wrkBusy_8 &&
	     wci_wciResponse_8$wget[33:32] != 2'd0 ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T ;

  // register wci_reqPend_9
  always@(MUX_wci_reqPend_9$write_1__SEL_1 or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_T_T or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T)
  begin
    case (1'b1) // synopsys parallel_case
      MUX_wci_reqPend_9$write_1__SEL_1: wci_reqPend_9$D_IN = 2'd0;
      WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_T_T:
	  wci_reqPend_9$D_IN = 2'd1;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T:
	  wci_reqPend_9$D_IN = 2'd2;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T:
	  wci_reqPend_9$D_IN = 2'd3;
      default: wci_reqPend_9$D_IN = 2'b10 /* unspecified value */ ;
    endcase
  end
  assign wci_reqPend_9$EN =
	     WILL_FIRE_RL_wci_wrkBusy_9 &&
	     wci_wciResponse_9$wget[33:32] != 2'd0 ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T ;

  // register wci_reqTO
  assign wci_reqTO$D_IN =
	     MUX_wci_reqTO$write_1__SEL_1 ?
	       MUX_wci_reqTO$write_1__VAL_1 :
	       3'd0 ;
  assign wci_reqTO$EN =
	     WILL_FIRE_RL_wci_wrkBusy &&
	     wci_wciResponse_wget__23_BITS_33_TO_32_24_EQ_0_ETC___d252 ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_T_F_F_T_T_T ;

  // register wci_reqTO_1
  assign wci_reqTO_1$D_IN =
	     MUX_wci_reqTO_1$write_1__SEL_1 ?
	       MUX_wci_reqTO_1$write_1__VAL_1 :
	       3'd0 ;
  assign wci_reqTO_1$EN =
	     WILL_FIRE_RL_wci_wrkBusy_1 &&
	     wci_wciResponse_1_wget__63_BITS_33_TO_32_64_EQ_ETC___d392 ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_T_F_F_T_T_T ;

  // register wci_reqTO_10
  assign wci_reqTO_10$D_IN =
	     MUX_wci_reqTO_10$write_1__SEL_1 ?
	       MUX_wci_reqTO_10$write_1__VAL_1 :
	       3'd0 ;
  assign wci_reqTO_10$EN =
	     WILL_FIRE_RL_wci_wrkBusy_10 &&
	     wci_wciResponse_10_wget__623_BITS_33_TO_32_624_ETC___d1652 ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T ;

  // register wci_reqTO_11
  assign wci_reqTO_11$D_IN =
	     MUX_wci_reqTO_11$write_1__SEL_1 ?
	       MUX_wci_reqTO_11$write_1__VAL_1 :
	       3'd0 ;
  assign wci_reqTO_11$EN =
	     WILL_FIRE_RL_wci_wrkBusy_11 &&
	     wci_wciResponse_11_wget__763_BITS_33_TO_32_764_ETC___d1792 ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T ;

  // register wci_reqTO_12
  assign wci_reqTO_12$D_IN =
	     MUX_wci_reqTO_12$write_1__SEL_1 ?
	       MUX_wci_reqTO_12$write_1__VAL_1 :
	       3'd0 ;
  assign wci_reqTO_12$EN =
	     WILL_FIRE_RL_wci_wrkBusy_12 &&
	     wci_wciResponse_12_wget__903_BITS_33_TO_32_904_ETC___d1932 ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T ;

  // register wci_reqTO_13
  assign wci_reqTO_13$D_IN =
	     MUX_wci_reqTO_13$write_1__SEL_1 ?
	       MUX_wci_reqTO_13$write_1__VAL_1 :
	       3'd0 ;
  assign wci_reqTO_13$EN =
	     WILL_FIRE_RL_wci_wrkBusy_13 &&
	     wci_wciResponse_13_wget__043_BITS_33_TO_32_044_ETC___d2072 ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T ;

  // register wci_reqTO_14
  assign wci_reqTO_14$D_IN =
	     MUX_wci_reqTO_14$write_1__SEL_1 ?
	       MUX_wci_reqTO_14$write_1__VAL_1 :
	       3'd0 ;
  assign wci_reqTO_14$EN =
	     WILL_FIRE_RL_wci_wrkBusy_14 &&
	     wci_wciResponse_14_wget__183_BITS_33_TO_32_184_ETC___d2212 ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T ;

  // register wci_reqTO_2
  assign wci_reqTO_2$D_IN =
	     MUX_wci_reqTO_2$write_1__SEL_1 ?
	       MUX_wci_reqTO_2$write_1__VAL_1 :
	       3'd0 ;
  assign wci_reqTO_2$EN =
	     WILL_FIRE_RL_wci_wrkBusy_2 &&
	     wci_wciResponse_2_wget__03_BITS_33_TO_32_04_EQ_ETC___d532 ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_F_F_T_T_T ;

  // register wci_reqTO_3
  assign wci_reqTO_3$D_IN =
	     MUX_wci_reqTO_3$write_1__SEL_1 ?
	       MUX_wci_reqTO_3$write_1__VAL_1 :
	       3'd0 ;
  assign wci_reqTO_3$EN =
	     WILL_FIRE_RL_wci_wrkBusy_3 &&
	     wci_wciResponse_3_wget__43_BITS_33_TO_32_44_EQ_ETC___d672 ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_F_F_T_T_T ;

  // register wci_reqTO_4
  assign wci_reqTO_4$D_IN =
	     MUX_wci_reqTO_4$write_1__SEL_1 ?
	       MUX_wci_reqTO_4$write_1__VAL_1 :
	       3'd0 ;
  assign wci_reqTO_4$EN =
	     WILL_FIRE_RL_wci_wrkBusy_4 &&
	     wci_wciResponse_4_wget__83_BITS_33_TO_32_84_EQ_ETC___d812 ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_F_F_T_T_T ;

  // register wci_reqTO_5
  assign wci_reqTO_5$D_IN =
	     MUX_wci_reqTO_5$write_1__SEL_1 ?
	       MUX_wci_reqTO_5$write_1__VAL_1 :
	       3'd0 ;
  assign wci_reqTO_5$EN =
	     WILL_FIRE_RL_wci_wrkBusy_5 &&
	     wci_wciResponse_5_wget__23_BITS_33_TO_32_24_EQ_ETC___d952 ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_F_T_T_T ;

  // register wci_reqTO_6
  assign wci_reqTO_6$D_IN =
	     MUX_wci_reqTO_6$write_1__SEL_1 ?
	       MUX_wci_reqTO_6$write_1__VAL_1 :
	       3'd0 ;
  assign wci_reqTO_6$EN =
	     WILL_FIRE_RL_wci_wrkBusy_6 &&
	     wci_wciResponse_6_wget__063_BITS_33_TO_32_064__ETC___d1092 ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_F_T_T_T ;

  // register wci_reqTO_7
  assign wci_reqTO_7$D_IN =
	     MUX_wci_reqTO_7$write_1__SEL_1 ?
	       MUX_wci_reqTO_7$write_1__VAL_1 :
	       3'd0 ;
  assign wci_reqTO_7$EN =
	     WILL_FIRE_RL_wci_wrkBusy_7 &&
	     wci_wciResponse_7_wget__203_BITS_33_TO_32_204__ETC___d1232 ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_F_T_T_T ;

  // register wci_reqTO_8
  assign wci_reqTO_8$D_IN =
	     MUX_wci_reqTO_8$write_1__SEL_1 ?
	       MUX_wci_reqTO_8$write_1__VAL_1 :
	       3'd0 ;
  assign wci_reqTO_8$EN =
	     WILL_FIRE_RL_wci_wrkBusy_8 &&
	     wci_wciResponse_8_wget__343_BITS_33_TO_32_344__ETC___d1372 ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_F_T_T_T ;

  // register wci_reqTO_9
  assign wci_reqTO_9$D_IN =
	     MUX_wci_reqTO_9$write_1__SEL_1 ?
	       MUX_wci_reqTO_9$write_1__VAL_1 :
	       3'd0 ;
  assign wci_reqTO_9$EN =
	     WILL_FIRE_RL_wci_wrkBusy_9 &&
	     wci_wciResponse_9_wget__483_BITS_33_TO_32_484__ETC___d1512 ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T ;

  // register wci_respTimr
  assign wci_respTimr$D_IN =
	     wci_reqF_c_r ? 32'd0 : MUX_wci_respTimr$write_1__VAL_2 ;
  assign wci_respTimr$EN = WILL_FIRE_RL_wci_wrkBusy || wci_reqF_c_r ;

  // register wci_respTimrAct
  assign wci_respTimrAct$D_IN = wci_reqF_c_r ;
  assign wci_respTimrAct$EN =
	     WILL_FIRE_RL_wci_wrkBusy &&
	     (!wci_respTimr_28_ULT_1_SL_wci_wTimeout_29_30___d5879 ||
	      wci_wciResponse$wget[33:32] != 2'd0) ||
	     wci_reqF_c_r ;

  // register wci_respTimrAct_1
  assign wci_respTimrAct_1$D_IN = wci_reqF_1_c_r ;
  assign wci_respTimrAct_1$EN =
	     WILL_FIRE_RL_wci_wrkBusy_1 &&
	     (!wci_respTimr_1_68_ULT_1_SL_wci_wTimeout_1_69_70___d5880 ||
	      wci_wciResponse_1$wget[33:32] != 2'd0) ||
	     wci_reqF_1_c_r ;

  // register wci_respTimrAct_10
  assign wci_respTimrAct_10$D_IN = wci_reqF_10_c_r ;
  assign wci_respTimrAct_10$EN =
	     WILL_FIRE_RL_wci_wrkBusy_10 &&
	     (!wci_respTimr_10_628_ULT_1_SL_wci_wTimeout_10_6_ETC___d5889 ||
	      wci_wciResponse_10$wget[33:32] != 2'd0) ||
	     wci_reqF_10_c_r ;

  // register wci_respTimrAct_11
  assign wci_respTimrAct_11$D_IN = wci_reqF_11_c_r ;
  assign wci_respTimrAct_11$EN =
	     WILL_FIRE_RL_wci_wrkBusy_11 &&
	     (!wci_respTimr_11_768_ULT_1_SL_wci_wTimeout_11_7_ETC___d5890 ||
	      wci_wciResponse_11$wget[33:32] != 2'd0) ||
	     wci_reqF_11_c_r ;

  // register wci_respTimrAct_12
  assign wci_respTimrAct_12$D_IN = wci_reqF_12_c_r ;
  assign wci_respTimrAct_12$EN =
	     WILL_FIRE_RL_wci_wrkBusy_12 &&
	     (!wci_respTimr_12_908_ULT_1_SL_wci_wTimeout_12_9_ETC___d5891 ||
	      wci_wciResponse_12$wget[33:32] != 2'd0) ||
	     wci_reqF_12_c_r ;

  // register wci_respTimrAct_13
  assign wci_respTimrAct_13$D_IN = wci_reqF_13_c_r ;
  assign wci_respTimrAct_13$EN =
	     WILL_FIRE_RL_wci_wrkBusy_13 &&
	     (!wci_respTimr_13_048_ULT_1_SL_wci_wTimeout_13_0_ETC___d5892 ||
	      wci_wciResponse_13$wget[33:32] != 2'd0) ||
	     wci_reqF_13_c_r ;

  // register wci_respTimrAct_14
  assign wci_respTimrAct_14$D_IN = wci_reqF_14_c_r ;
  assign wci_respTimrAct_14$EN =
	     WILL_FIRE_RL_wci_wrkBusy_14 &&
	     (!wci_respTimr_14_188_ULT_1_SL_wci_wTimeout_14_1_ETC___d5893 ||
	      wci_wciResponse_14$wget[33:32] != 2'd0) ||
	     wci_reqF_14_c_r ;

  // register wci_respTimrAct_2
  assign wci_respTimrAct_2$D_IN = wci_reqF_2_c_r ;
  assign wci_respTimrAct_2$EN =
	     WILL_FIRE_RL_wci_wrkBusy_2 &&
	     (!wci_respTimr_2_08_ULT_1_SL_wci_wTimeout_2_09_10___d5881 ||
	      wci_wciResponse_2$wget[33:32] != 2'd0) ||
	     wci_reqF_2_c_r ;

  // register wci_respTimrAct_3
  assign wci_respTimrAct_3$D_IN = wci_reqF_3_c_r ;
  assign wci_respTimrAct_3$EN =
	     WILL_FIRE_RL_wci_wrkBusy_3 &&
	     (!wci_respTimr_3_48_ULT_1_SL_wci_wTimeout_3_49_50___d5882 ||
	      wci_wciResponse_3$wget[33:32] != 2'd0) ||
	     wci_reqF_3_c_r ;

  // register wci_respTimrAct_4
  assign wci_respTimrAct_4$D_IN = wci_reqF_4_c_r ;
  assign wci_respTimrAct_4$EN =
	     WILL_FIRE_RL_wci_wrkBusy_4 &&
	     (!wci_respTimr_4_88_ULT_1_SL_wci_wTimeout_4_89_90___d5883 ||
	      wci_wciResponse_4$wget[33:32] != 2'd0) ||
	     wci_reqF_4_c_r ;

  // register wci_respTimrAct_5
  assign wci_respTimrAct_5$D_IN = wci_reqF_5_c_r ;
  assign wci_respTimrAct_5$EN =
	     WILL_FIRE_RL_wci_wrkBusy_5 &&
	     (!wci_respTimr_5_28_ULT_1_SL_wci_wTimeout_5_29_30___d5884 ||
	      wci_wciResponse_5$wget[33:32] != 2'd0) ||
	     wci_reqF_5_c_r ;

  // register wci_respTimrAct_6
  assign wci_respTimrAct_6$D_IN = wci_reqF_6_c_r ;
  assign wci_respTimrAct_6$EN =
	     WILL_FIRE_RL_wci_wrkBusy_6 &&
	     (!wci_respTimr_6_068_ULT_1_SL_wci_wTimeout_6_069_ETC___d5885 ||
	      wci_wciResponse_6$wget[33:32] != 2'd0) ||
	     wci_reqF_6_c_r ;

  // register wci_respTimrAct_7
  assign wci_respTimrAct_7$D_IN = wci_reqF_7_c_r ;
  assign wci_respTimrAct_7$EN =
	     WILL_FIRE_RL_wci_wrkBusy_7 &&
	     (!wci_respTimr_7_208_ULT_1_SL_wci_wTimeout_7_209_ETC___d5886 ||
	      wci_wciResponse_7$wget[33:32] != 2'd0) ||
	     wci_reqF_7_c_r ;

  // register wci_respTimrAct_8
  assign wci_respTimrAct_8$D_IN = wci_reqF_8_c_r ;
  assign wci_respTimrAct_8$EN =
	     WILL_FIRE_RL_wci_wrkBusy_8 &&
	     (!wci_respTimr_8_348_ULT_1_SL_wci_wTimeout_8_349_ETC___d5887 ||
	      wci_wciResponse_8$wget[33:32] != 2'd0) ||
	     wci_reqF_8_c_r ;

  // register wci_respTimrAct_9
  assign wci_respTimrAct_9$D_IN = wci_reqF_9_c_r ;
  assign wci_respTimrAct_9$EN =
	     WILL_FIRE_RL_wci_wrkBusy_9 &&
	     (!wci_respTimr_9_488_ULT_1_SL_wci_wTimeout_9_489_ETC___d5888 ||
	      wci_wciResponse_9$wget[33:32] != 2'd0) ||
	     wci_reqF_9_c_r ;

  // register wci_respTimr_1
  assign wci_respTimr_1$D_IN =
	     wci_reqF_1_c_r ? 32'd0 : MUX_wci_respTimr_1$write_1__VAL_2 ;
  assign wci_respTimr_1$EN = WILL_FIRE_RL_wci_wrkBusy_1 || wci_reqF_1_c_r ;

  // register wci_respTimr_10
  assign wci_respTimr_10$D_IN =
	     wci_reqF_10_c_r ? 32'd0 : MUX_wci_respTimr_10$write_1__VAL_2 ;
  assign wci_respTimr_10$EN = WILL_FIRE_RL_wci_wrkBusy_10 || wci_reqF_10_c_r ;

  // register wci_respTimr_11
  assign wci_respTimr_11$D_IN =
	     wci_reqF_11_c_r ? 32'd0 : MUX_wci_respTimr_11$write_1__VAL_2 ;
  assign wci_respTimr_11$EN = WILL_FIRE_RL_wci_wrkBusy_11 || wci_reqF_11_c_r ;

  // register wci_respTimr_12
  assign wci_respTimr_12$D_IN =
	     wci_reqF_12_c_r ? 32'd0 : MUX_wci_respTimr_12$write_1__VAL_2 ;
  assign wci_respTimr_12$EN = WILL_FIRE_RL_wci_wrkBusy_12 || wci_reqF_12_c_r ;

  // register wci_respTimr_13
  assign wci_respTimr_13$D_IN =
	     wci_reqF_13_c_r ? 32'd0 : MUX_wci_respTimr_13$write_1__VAL_2 ;
  assign wci_respTimr_13$EN = WILL_FIRE_RL_wci_wrkBusy_13 || wci_reqF_13_c_r ;

  // register wci_respTimr_14
  assign wci_respTimr_14$D_IN =
	     wci_reqF_14_c_r ? 32'd0 : MUX_wci_respTimr_14$write_1__VAL_2 ;
  assign wci_respTimr_14$EN = WILL_FIRE_RL_wci_wrkBusy_14 || wci_reqF_14_c_r ;

  // register wci_respTimr_2
  assign wci_respTimr_2$D_IN =
	     wci_reqF_2_c_r ? 32'd0 : MUX_wci_respTimr_2$write_1__VAL_2 ;
  assign wci_respTimr_2$EN = WILL_FIRE_RL_wci_wrkBusy_2 || wci_reqF_2_c_r ;

  // register wci_respTimr_3
  assign wci_respTimr_3$D_IN =
	     wci_reqF_3_c_r ? 32'd0 : MUX_wci_respTimr_3$write_1__VAL_2 ;
  assign wci_respTimr_3$EN = WILL_FIRE_RL_wci_wrkBusy_3 || wci_reqF_3_c_r ;

  // register wci_respTimr_4
  assign wci_respTimr_4$D_IN =
	     wci_reqF_4_c_r ? 32'd0 : MUX_wci_respTimr_4$write_1__VAL_2 ;
  assign wci_respTimr_4$EN = WILL_FIRE_RL_wci_wrkBusy_4 || wci_reqF_4_c_r ;

  // register wci_respTimr_5
  assign wci_respTimr_5$D_IN =
	     wci_reqF_5_c_r ? 32'd0 : MUX_wci_respTimr_5$write_1__VAL_2 ;
  assign wci_respTimr_5$EN = WILL_FIRE_RL_wci_wrkBusy_5 || wci_reqF_5_c_r ;

  // register wci_respTimr_6
  assign wci_respTimr_6$D_IN =
	     wci_reqF_6_c_r ? 32'd0 : MUX_wci_respTimr_6$write_1__VAL_2 ;
  assign wci_respTimr_6$EN = WILL_FIRE_RL_wci_wrkBusy_6 || wci_reqF_6_c_r ;

  // register wci_respTimr_7
  assign wci_respTimr_7$D_IN =
	     wci_reqF_7_c_r ? 32'd0 : MUX_wci_respTimr_7$write_1__VAL_2 ;
  assign wci_respTimr_7$EN = WILL_FIRE_RL_wci_wrkBusy_7 || wci_reqF_7_c_r ;

  // register wci_respTimr_8
  assign wci_respTimr_8$D_IN =
	     wci_reqF_8_c_r ? 32'd0 : MUX_wci_respTimr_8$write_1__VAL_2 ;
  assign wci_respTimr_8$EN = WILL_FIRE_RL_wci_wrkBusy_8 || wci_reqF_8_c_r ;

  // register wci_respTimr_9
  assign wci_respTimr_9$D_IN =
	     wci_reqF_9_c_r ? 32'd0 : MUX_wci_respTimr_9$write_1__VAL_2 ;
  assign wci_respTimr_9$EN = WILL_FIRE_RL_wci_wrkBusy_9 || wci_reqF_9_c_r ;

  // register wci_sThreadBusy_d
  assign wci_sThreadBusy_d$D_IN = wci_Vm_0_SThreadBusy ;
  assign wci_sThreadBusy_d$EN = 1'd1 ;

  // register wci_sThreadBusy_d_1
  assign wci_sThreadBusy_d_1$D_IN = wci_Vm_1_SThreadBusy ;
  assign wci_sThreadBusy_d_1$EN = 1'd1 ;

  // register wci_sThreadBusy_d_10
  assign wci_sThreadBusy_d_10$D_IN = wci_Vm_10_SThreadBusy ;
  assign wci_sThreadBusy_d_10$EN = 1'd1 ;

  // register wci_sThreadBusy_d_11
  assign wci_sThreadBusy_d_11$D_IN = wci_Vm_11_SThreadBusy ;
  assign wci_sThreadBusy_d_11$EN = 1'd1 ;

  // register wci_sThreadBusy_d_12
  assign wci_sThreadBusy_d_12$D_IN = wci_Vm_12_SThreadBusy ;
  assign wci_sThreadBusy_d_12$EN = 1'd1 ;

  // register wci_sThreadBusy_d_13
  assign wci_sThreadBusy_d_13$D_IN = wci_Vm_13_SThreadBusy ;
  assign wci_sThreadBusy_d_13$EN = 1'd1 ;

  // register wci_sThreadBusy_d_14
  assign wci_sThreadBusy_d_14$D_IN = wci_Vm_14_SThreadBusy ;
  assign wci_sThreadBusy_d_14$EN = 1'd1 ;

  // register wci_sThreadBusy_d_2
  assign wci_sThreadBusy_d_2$D_IN = wci_Vm_2_SThreadBusy ;
  assign wci_sThreadBusy_d_2$EN = 1'd1 ;

  // register wci_sThreadBusy_d_3
  assign wci_sThreadBusy_d_3$D_IN = wci_Vm_3_SThreadBusy ;
  assign wci_sThreadBusy_d_3$EN = 1'd1 ;

  // register wci_sThreadBusy_d_4
  assign wci_sThreadBusy_d_4$D_IN = wci_Vm_4_SThreadBusy ;
  assign wci_sThreadBusy_d_4$EN = 1'd1 ;

  // register wci_sThreadBusy_d_5
  assign wci_sThreadBusy_d_5$D_IN = wci_Vm_5_SThreadBusy ;
  assign wci_sThreadBusy_d_5$EN = 1'd1 ;

  // register wci_sThreadBusy_d_6
  assign wci_sThreadBusy_d_6$D_IN = wci_Vm_6_SThreadBusy ;
  assign wci_sThreadBusy_d_6$EN = 1'd1 ;

  // register wci_sThreadBusy_d_7
  assign wci_sThreadBusy_d_7$D_IN = wci_Vm_7_SThreadBusy ;
  assign wci_sThreadBusy_d_7$EN = 1'd1 ;

  // register wci_sThreadBusy_d_8
  assign wci_sThreadBusy_d_8$D_IN = wci_Vm_8_SThreadBusy ;
  assign wci_sThreadBusy_d_8$EN = 1'd1 ;

  // register wci_sThreadBusy_d_9
  assign wci_sThreadBusy_d_9$D_IN = wci_Vm_9_SThreadBusy ;
  assign wci_sThreadBusy_d_9$EN = 1'd1 ;

  // register wci_sfCap
  assign wci_sfCap$D_IN = wci_sfCapSet ;
  assign wci_sfCap$EN = wci_sfCapSet || wci_sfCapClear ;

  // register wci_sfCapClear
  assign wci_sfCapClear$D_IN = wci_sfCapClear_1$whas ;
  assign wci_sfCapClear$EN = 1'd1 ;

  // register wci_sfCapClear_10
  assign wci_sfCapClear_10$D_IN = wci_sfCapClear_10_1$whas ;
  assign wci_sfCapClear_10$EN = 1'd1 ;

  // register wci_sfCapClear_11
  assign wci_sfCapClear_11$D_IN = wci_sfCapClear_11_1$whas ;
  assign wci_sfCapClear_11$EN = 1'd1 ;

  // register wci_sfCapClear_12
  assign wci_sfCapClear_12$D_IN = wci_sfCapClear_12_1$whas ;
  assign wci_sfCapClear_12$EN = 1'd1 ;

  // register wci_sfCapClear_13
  assign wci_sfCapClear_13$D_IN = wci_sfCapClear_13_1$whas ;
  assign wci_sfCapClear_13$EN = 1'd1 ;

  // register wci_sfCapClear_14
  assign wci_sfCapClear_14$D_IN = wci_sfCapClear_14_1$whas ;
  assign wci_sfCapClear_14$EN = 1'd1 ;

  // register wci_sfCapClear_1_1
  assign wci_sfCapClear_1_1$D_IN = wci_sfCapClear_1_2$whas ;
  assign wci_sfCapClear_1_1$EN = 1'd1 ;

  // register wci_sfCapClear_2
  assign wci_sfCapClear_2$D_IN = wci_sfCapClear_2_1$whas ;
  assign wci_sfCapClear_2$EN = 1'd1 ;

  // register wci_sfCapClear_3
  assign wci_sfCapClear_3$D_IN = wci_sfCapClear_3_1$whas ;
  assign wci_sfCapClear_3$EN = 1'd1 ;

  // register wci_sfCapClear_4
  assign wci_sfCapClear_4$D_IN = wci_sfCapClear_4_1$whas ;
  assign wci_sfCapClear_4$EN = 1'd1 ;

  // register wci_sfCapClear_5
  assign wci_sfCapClear_5$D_IN = wci_sfCapClear_5_1$whas ;
  assign wci_sfCapClear_5$EN = 1'd1 ;

  // register wci_sfCapClear_6
  assign wci_sfCapClear_6$D_IN = wci_sfCapClear_6_1$whas ;
  assign wci_sfCapClear_6$EN = 1'd1 ;

  // register wci_sfCapClear_7
  assign wci_sfCapClear_7$D_IN = wci_sfCapClear_7_1$whas ;
  assign wci_sfCapClear_7$EN = 1'd1 ;

  // register wci_sfCapClear_8
  assign wci_sfCapClear_8$D_IN = wci_sfCapClear_8_1$whas ;
  assign wci_sfCapClear_8$EN = 1'd1 ;

  // register wci_sfCapClear_9
  assign wci_sfCapClear_9$D_IN = wci_sfCapClear_9_1$whas ;
  assign wci_sfCapClear_9$EN = 1'd1 ;

  // register wci_sfCapSet
  assign wci_sfCapSet$D_IN = wci_Vm_0_SFlag[0] ;
  assign wci_sfCapSet$EN = 1'd1 ;

  // register wci_sfCapSet_10
  assign wci_sfCapSet_10$D_IN = wci_Vm_10_SFlag[0] ;
  assign wci_sfCapSet_10$EN = 1'd1 ;

  // register wci_sfCapSet_11
  assign wci_sfCapSet_11$D_IN = wci_Vm_11_SFlag[0] ;
  assign wci_sfCapSet_11$EN = 1'd1 ;

  // register wci_sfCapSet_12
  assign wci_sfCapSet_12$D_IN = wci_Vm_12_SFlag[0] ;
  assign wci_sfCapSet_12$EN = 1'd1 ;

  // register wci_sfCapSet_13
  assign wci_sfCapSet_13$D_IN = wci_Vm_13_SFlag[0] ;
  assign wci_sfCapSet_13$EN = 1'd1 ;

  // register wci_sfCapSet_14
  assign wci_sfCapSet_14$D_IN = wci_Vm_14_SFlag[0] ;
  assign wci_sfCapSet_14$EN = 1'd1 ;

  // register wci_sfCapSet_1_1
  assign wci_sfCapSet_1_1$D_IN = wci_Vm_1_SFlag[0] ;
  assign wci_sfCapSet_1_1$EN = 1'd1 ;

  // register wci_sfCapSet_2
  assign wci_sfCapSet_2$D_IN = wci_Vm_2_SFlag[0] ;
  assign wci_sfCapSet_2$EN = 1'd1 ;

  // register wci_sfCapSet_3
  assign wci_sfCapSet_3$D_IN = wci_Vm_3_SFlag[0] ;
  assign wci_sfCapSet_3$EN = 1'd1 ;

  // register wci_sfCapSet_4
  assign wci_sfCapSet_4$D_IN = wci_Vm_4_SFlag[0] ;
  assign wci_sfCapSet_4$EN = 1'd1 ;

  // register wci_sfCapSet_5
  assign wci_sfCapSet_5$D_IN = wci_Vm_5_SFlag[0] ;
  assign wci_sfCapSet_5$EN = 1'd1 ;

  // register wci_sfCapSet_6
  assign wci_sfCapSet_6$D_IN = wci_Vm_6_SFlag[0] ;
  assign wci_sfCapSet_6$EN = 1'd1 ;

  // register wci_sfCapSet_7
  assign wci_sfCapSet_7$D_IN = wci_Vm_7_SFlag[0] ;
  assign wci_sfCapSet_7$EN = 1'd1 ;

  // register wci_sfCapSet_8
  assign wci_sfCapSet_8$D_IN = wci_Vm_8_SFlag[0] ;
  assign wci_sfCapSet_8$EN = 1'd1 ;

  // register wci_sfCapSet_9
  assign wci_sfCapSet_9$D_IN = wci_Vm_9_SFlag[0] ;
  assign wci_sfCapSet_9$EN = 1'd1 ;

  // register wci_sfCap_1
  assign wci_sfCap_1$D_IN = wci_sfCapSet_1_1 ;
  assign wci_sfCap_1$EN = wci_sfCapSet_1_1 || wci_sfCapClear_1_1 ;

  // register wci_sfCap_10
  assign wci_sfCap_10$D_IN = wci_sfCapSet_10 ;
  assign wci_sfCap_10$EN = wci_sfCapSet_10 || wci_sfCapClear_10 ;

  // register wci_sfCap_11
  assign wci_sfCap_11$D_IN = wci_sfCapSet_11 ;
  assign wci_sfCap_11$EN = wci_sfCapSet_11 || wci_sfCapClear_11 ;

  // register wci_sfCap_12
  assign wci_sfCap_12$D_IN = wci_sfCapSet_12 ;
  assign wci_sfCap_12$EN = wci_sfCapSet_12 || wci_sfCapClear_12 ;

  // register wci_sfCap_13
  assign wci_sfCap_13$D_IN = wci_sfCapSet_13 ;
  assign wci_sfCap_13$EN = wci_sfCapSet_13 || wci_sfCapClear_13 ;

  // register wci_sfCap_14
  assign wci_sfCap_14$D_IN = wci_sfCapSet_14 ;
  assign wci_sfCap_14$EN = wci_sfCapSet_14 || wci_sfCapClear_14 ;

  // register wci_sfCap_2
  assign wci_sfCap_2$D_IN = wci_sfCapSet_2 ;
  assign wci_sfCap_2$EN = wci_sfCapSet_2 || wci_sfCapClear_2 ;

  // register wci_sfCap_3
  assign wci_sfCap_3$D_IN = wci_sfCapSet_3 ;
  assign wci_sfCap_3$EN = wci_sfCapSet_3 || wci_sfCapClear_3 ;

  // register wci_sfCap_4
  assign wci_sfCap_4$D_IN = wci_sfCapSet_4 ;
  assign wci_sfCap_4$EN = wci_sfCapSet_4 || wci_sfCapClear_4 ;

  // register wci_sfCap_5
  assign wci_sfCap_5$D_IN = wci_sfCapSet_5 ;
  assign wci_sfCap_5$EN = wci_sfCapSet_5 || wci_sfCapClear_5 ;

  // register wci_sfCap_6
  assign wci_sfCap_6$D_IN = wci_sfCapSet_6 ;
  assign wci_sfCap_6$EN = wci_sfCapSet_6 || wci_sfCapClear_6 ;

  // register wci_sfCap_7
  assign wci_sfCap_7$D_IN = wci_sfCapSet_7 ;
  assign wci_sfCap_7$EN = wci_sfCapSet_7 || wci_sfCapClear_7 ;

  // register wci_sfCap_8
  assign wci_sfCap_8$D_IN = wci_sfCapSet_8 ;
  assign wci_sfCap_8$EN = wci_sfCapSet_8 || wci_sfCapClear_8 ;

  // register wci_sfCap_9
  assign wci_sfCap_9$D_IN = wci_sfCapSet_9 ;
  assign wci_sfCap_9$EN = wci_sfCapSet_9 || wci_sfCapClear_9 ;

  // register wci_slvPresent
  assign wci_slvPresent$D_IN = wci_Vm_0_SFlag[1] ;
  assign wci_slvPresent$EN = 1'd1 ;

  // register wci_slvPresent_1
  assign wci_slvPresent_1$D_IN = wci_Vm_1_SFlag[1] ;
  assign wci_slvPresent_1$EN = 1'd1 ;

  // register wci_slvPresent_10
  assign wci_slvPresent_10$D_IN = wci_Vm_10_SFlag[1] ;
  assign wci_slvPresent_10$EN = 1'd1 ;

  // register wci_slvPresent_11
  assign wci_slvPresent_11$D_IN = wci_Vm_11_SFlag[1] ;
  assign wci_slvPresent_11$EN = 1'd1 ;

  // register wci_slvPresent_12
  assign wci_slvPresent_12$D_IN = wci_Vm_12_SFlag[1] ;
  assign wci_slvPresent_12$EN = 1'd1 ;

  // register wci_slvPresent_13
  assign wci_slvPresent_13$D_IN = wci_Vm_13_SFlag[1] ;
  assign wci_slvPresent_13$EN = 1'd1 ;

  // register wci_slvPresent_14
  assign wci_slvPresent_14$D_IN = wci_Vm_14_SFlag[1] ;
  assign wci_slvPresent_14$EN = 1'd1 ;

  // register wci_slvPresent_2
  assign wci_slvPresent_2$D_IN = wci_Vm_2_SFlag[1] ;
  assign wci_slvPresent_2$EN = 1'd1 ;

  // register wci_slvPresent_3
  assign wci_slvPresent_3$D_IN = wci_Vm_3_SFlag[1] ;
  assign wci_slvPresent_3$EN = 1'd1 ;

  // register wci_slvPresent_4
  assign wci_slvPresent_4$D_IN = wci_Vm_4_SFlag[1] ;
  assign wci_slvPresent_4$EN = 1'd1 ;

  // register wci_slvPresent_5
  assign wci_slvPresent_5$D_IN = wci_Vm_5_SFlag[1] ;
  assign wci_slvPresent_5$EN = 1'd1 ;

  // register wci_slvPresent_6
  assign wci_slvPresent_6$D_IN = wci_Vm_6_SFlag[1] ;
  assign wci_slvPresent_6$EN = 1'd1 ;

  // register wci_slvPresent_7
  assign wci_slvPresent_7$D_IN = wci_Vm_7_SFlag[1] ;
  assign wci_slvPresent_7$EN = 1'd1 ;

  // register wci_slvPresent_8
  assign wci_slvPresent_8$D_IN = wci_Vm_8_SFlag[1] ;
  assign wci_slvPresent_8$EN = 1'd1 ;

  // register wci_slvPresent_9
  assign wci_slvPresent_9$D_IN = wci_Vm_9_SFlag[1] ;
  assign wci_slvPresent_9$EN = 1'd1 ;

  // register wci_wReset_n
  assign wci_wReset_n$D_IN = cpReq[59] ;
  assign wci_wReset_n$EN =
	     WILL_FIRE_RL_cpDispatch_F_F_T_T_F_F_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_T_F_F_T_T_T ;

  // register wci_wReset_n_1
  assign wci_wReset_n_1$D_IN = cpReq[59] ;
  assign wci_wReset_n_1$EN =
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_T_F_F_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_T_F_F_T_T_T ;

  // register wci_wReset_n_10
  assign wci_wReset_n_10$D_IN = cpReq[59] ;
  assign wci_wReset_n_10$EN =
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T ;

  // register wci_wReset_n_11
  assign wci_wReset_n_11$D_IN = cpReq[59] ;
  assign wci_wReset_n_11$EN =
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T ;

  // register wci_wReset_n_12
  assign wci_wReset_n_12$D_IN = cpReq[59] ;
  assign wci_wReset_n_12$EN =
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T ;

  // register wci_wReset_n_13
  assign wci_wReset_n_13$D_IN = cpReq[59] ;
  assign wci_wReset_n_13$EN =
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T ;

  // register wci_wReset_n_14
  assign wci_wReset_n_14$D_IN = cpReq[59] ;
  assign wci_wReset_n_14$EN =
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T ;

  // register wci_wReset_n_2
  assign wci_wReset_n_2$D_IN = cpReq[59] ;
  assign wci_wReset_n_2$EN =
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_F_F_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_F_F_T_T_T ;

  // register wci_wReset_n_3
  assign wci_wReset_n_3$D_IN = cpReq[59] ;
  assign wci_wReset_n_3$EN =
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_F_F_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_F_F_T_T_T ;

  // register wci_wReset_n_4
  assign wci_wReset_n_4$D_IN = cpReq[59] ;
  assign wci_wReset_n_4$EN =
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_F_F_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_F_F_T_T_T ;

  // register wci_wReset_n_5
  assign wci_wReset_n_5$D_IN = cpReq[59] ;
  assign wci_wReset_n_5$EN =
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_F_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_F_T_T_T ;

  // register wci_wReset_n_6
  assign wci_wReset_n_6$D_IN = cpReq[59] ;
  assign wci_wReset_n_6$EN =
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_F_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_F_T_T_T ;

  // register wci_wReset_n_7
  assign wci_wReset_n_7$D_IN = cpReq[59] ;
  assign wci_wReset_n_7$EN =
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_F_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_F_T_T_T ;

  // register wci_wReset_n_8
  assign wci_wReset_n_8$D_IN = cpReq[59] ;
  assign wci_wReset_n_8$EN =
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_F_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_F_T_T_T ;

  // register wci_wReset_n_9
  assign wci_wReset_n_9$D_IN = cpReq[59] ;
  assign wci_wReset_n_9$EN =
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_F_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T ;

  // register wci_wStatus
  assign wci_wStatus$D_IN =
	     { 4'b0,
	       !wci_lastOpWrite[1] || wci_lastOpWrite[0],
	       IF_wci_lastControlOp_13_BIT_3_14_THEN_wci_last_ETC___d328 } ;
  assign wci_wStatus$EN = 1'd1 ;

  // register wci_wStatus_1
  assign wci_wStatus_1$D_IN =
	     { 4'b0,
	       !wci_lastOpWrite_1[1] || wci_lastOpWrite_1[0],
	       IF_wci_lastControlOp_1_53_BIT_3_54_THEN_wci_la_ETC___d468 } ;
  assign wci_wStatus_1$EN = 1'd1 ;

  // register wci_wStatus_10
  assign wci_wStatus_10$D_IN =
	     { 4'b0,
	       !wci_lastOpWrite_10[1] || wci_lastOpWrite_10[0],
	       IF_wci_lastControlOp_10_713_BIT_3_714_THEN_wci_ETC___d1728 } ;
  assign wci_wStatus_10$EN = 1'd1 ;

  // register wci_wStatus_11
  assign wci_wStatus_11$D_IN =
	     { 4'b0,
	       !wci_lastOpWrite_11[1] || wci_lastOpWrite_11[0],
	       IF_wci_lastControlOp_11_853_BIT_3_854_THEN_wci_ETC___d1868 } ;
  assign wci_wStatus_11$EN = 1'd1 ;

  // register wci_wStatus_12
  assign wci_wStatus_12$D_IN =
	     { 4'b0,
	       !wci_lastOpWrite_12[1] || wci_lastOpWrite_12[0],
	       IF_wci_lastControlOp_12_993_BIT_3_994_THEN_wci_ETC___d2008 } ;
  assign wci_wStatus_12$EN = 1'd1 ;

  // register wci_wStatus_13
  assign wci_wStatus_13$D_IN =
	     { 4'b0,
	       !wci_lastOpWrite_13[1] || wci_lastOpWrite_13[0],
	       IF_wci_lastControlOp_13_133_BIT_3_134_THEN_wci_ETC___d2148 } ;
  assign wci_wStatus_13$EN = 1'd1 ;

  // register wci_wStatus_14
  assign wci_wStatus_14$D_IN =
	     { 4'b0,
	       !wci_lastOpWrite_14[1] || wci_lastOpWrite_14[0],
	       IF_wci_lastControlOp_14_273_BIT_3_274_THEN_wci_ETC___d2288 } ;
  assign wci_wStatus_14$EN = 1'd1 ;

  // register wci_wStatus_2
  assign wci_wStatus_2$D_IN =
	     { 4'b0,
	       !wci_lastOpWrite_2[1] || wci_lastOpWrite_2[0],
	       IF_wci_lastControlOp_2_93_BIT_3_94_THEN_wci_la_ETC___d608 } ;
  assign wci_wStatus_2$EN = 1'd1 ;

  // register wci_wStatus_3
  assign wci_wStatus_3$D_IN =
	     { 4'b0,
	       !wci_lastOpWrite_3[1] || wci_lastOpWrite_3[0],
	       IF_wci_lastControlOp_3_33_BIT_3_34_THEN_wci_la_ETC___d748 } ;
  assign wci_wStatus_3$EN = 1'd1 ;

  // register wci_wStatus_4
  assign wci_wStatus_4$D_IN =
	     { 4'b0,
	       !wci_lastOpWrite_4[1] || wci_lastOpWrite_4[0],
	       IF_wci_lastControlOp_4_73_BIT_3_74_THEN_wci_la_ETC___d888 } ;
  assign wci_wStatus_4$EN = 1'd1 ;

  // register wci_wStatus_5
  assign wci_wStatus_5$D_IN =
	     { 4'b0,
	       !wci_lastOpWrite_5[1] || wci_lastOpWrite_5[0],
	       IF_wci_lastControlOp_5_013_BIT_3_014_THEN_wci__ETC___d1028 } ;
  assign wci_wStatus_5$EN = 1'd1 ;

  // register wci_wStatus_6
  assign wci_wStatus_6$D_IN =
	     { 4'b0,
	       !wci_lastOpWrite_6[1] || wci_lastOpWrite_6[0],
	       IF_wci_lastControlOp_6_153_BIT_3_154_THEN_wci__ETC___d1168 } ;
  assign wci_wStatus_6$EN = 1'd1 ;

  // register wci_wStatus_7
  assign wci_wStatus_7$D_IN =
	     { 4'b0,
	       !wci_lastOpWrite_7[1] || wci_lastOpWrite_7[0],
	       IF_wci_lastControlOp_7_293_BIT_3_294_THEN_wci__ETC___d1308 } ;
  assign wci_wStatus_7$EN = 1'd1 ;

  // register wci_wStatus_8
  assign wci_wStatus_8$D_IN =
	     { 4'b0,
	       !wci_lastOpWrite_8[1] || wci_lastOpWrite_8[0],
	       IF_wci_lastControlOp_8_433_BIT_3_434_THEN_wci__ETC___d1448 } ;
  assign wci_wStatus_8$EN = 1'd1 ;

  // register wci_wStatus_9
  assign wci_wStatus_9$D_IN =
	     { 4'b0,
	       !wci_lastOpWrite_9[1] || wci_lastOpWrite_9[0],
	       IF_wci_lastControlOp_9_573_BIT_3_574_THEN_wci__ETC___d1588 } ;
  assign wci_wStatus_9$EN = 1'd1 ;

  // register wci_wTimeout
  assign wci_wTimeout$D_IN = cpReq[32:28] ;
  assign wci_wTimeout$EN =
	     WILL_FIRE_RL_cpDispatch_F_F_T_T_F_F_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_T_F_F_T_T_T ;

  // register wci_wTimeout_1
  assign wci_wTimeout_1$D_IN = cpReq[32:28] ;
  assign wci_wTimeout_1$EN =
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_T_F_F_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_T_F_F_T_T_T ;

  // register wci_wTimeout_10
  assign wci_wTimeout_10$D_IN = cpReq[32:28] ;
  assign wci_wTimeout_10$EN =
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T ;

  // register wci_wTimeout_11
  assign wci_wTimeout_11$D_IN = cpReq[32:28] ;
  assign wci_wTimeout_11$EN =
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T ;

  // register wci_wTimeout_12
  assign wci_wTimeout_12$D_IN = cpReq[32:28] ;
  assign wci_wTimeout_12$EN =
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T ;

  // register wci_wTimeout_13
  assign wci_wTimeout_13$D_IN = cpReq[32:28] ;
  assign wci_wTimeout_13$EN =
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T ;

  // register wci_wTimeout_14
  assign wci_wTimeout_14$D_IN = cpReq[32:28] ;
  assign wci_wTimeout_14$EN =
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T ;

  // register wci_wTimeout_2
  assign wci_wTimeout_2$D_IN = cpReq[32:28] ;
  assign wci_wTimeout_2$EN =
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_F_F_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_F_F_T_T_T ;

  // register wci_wTimeout_3
  assign wci_wTimeout_3$D_IN = cpReq[32:28] ;
  assign wci_wTimeout_3$EN =
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_F_F_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_F_F_T_T_T ;

  // register wci_wTimeout_4
  assign wci_wTimeout_4$D_IN = cpReq[32:28] ;
  assign wci_wTimeout_4$EN =
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_F_F_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_F_F_T_T_T ;

  // register wci_wTimeout_5
  assign wci_wTimeout_5$D_IN = cpReq[32:28] ;
  assign wci_wTimeout_5$EN =
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_F_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_F_T_T_T ;

  // register wci_wTimeout_6
  assign wci_wTimeout_6$D_IN = cpReq[32:28] ;
  assign wci_wTimeout_6$EN =
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_F_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_F_T_T_T ;

  // register wci_wTimeout_7
  assign wci_wTimeout_7$D_IN = cpReq[32:28] ;
  assign wci_wTimeout_7$EN =
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_F_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_F_T_T_T ;

  // register wci_wTimeout_8
  assign wci_wTimeout_8$D_IN = cpReq[32:28] ;
  assign wci_wTimeout_8$EN =
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_F_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_F_T_T_T ;

  // register wci_wTimeout_9
  assign wci_wTimeout_9$D_IN = cpReq[32:28] ;
  assign wci_wTimeout_9$EN =
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_F_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T ;

  // register wrkAct
  always@(MUX_wrkAct$write_1__SEL_1 or
	  _theResult_____1__h76796 or
	  MUX_wrkAct$write_1__SEL_2 or
	  _theResult_____1__h76814 or MUX_wrkAct$write_1__SEL_3)
  begin
    case (1'b1) // synopsys parallel_case
      MUX_wrkAct$write_1__SEL_1: wrkAct$D_IN = _theResult_____1__h76796;
      MUX_wrkAct$write_1__SEL_2: wrkAct$D_IN = _theResult_____1__h76814;
      MUX_wrkAct$write_1__SEL_3: wrkAct$D_IN = 4'd0;
      default: wrkAct$D_IN = 4'b1010 /* unspecified value */ ;
    endcase
  end
  assign wrkAct$EN =
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_F_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_F_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_F_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_F_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_F_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_F_F_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_F_F_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_F_F_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_T_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_T_F_F_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_T_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_T_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_T_F_F_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_T_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_F_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_F_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_F_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_F_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_F_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_F_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_F_F_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_F_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_F_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_F_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_F_F_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_F_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_F_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_F_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_F_F_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_F_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_F_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_F_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_T_F_F_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_T_F_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_T_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_T_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_T_F_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_T_F_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_T_T_T ||
	     WILL_FIRE_RL_completeWorkerRead ||
	     WILL_FIRE_RL_completeWorkerWrite ;

  // submodule adminResp1F
  assign adminResp1F$D_IN =
	     { cpReq[11:4] == 8'h0 || cpReq[11:4] == 8'h04 ||
	       cpReq[11:4] == 8'h08 ||
	       cpReq[11:4] == 8'h0C ||
	       cpReq[11:4] == 8'h10 ||
	       cpReq[11:4] == 8'h14 ||
	       cpReq[11:4] == 8'h18 ||
	       cpReq[11:4] == 8'h1C ||
	       cpReq[11:4] == 8'h20 ||
	       cpReq[11:4] == 8'h24 ||
	       cpReq[11:4] == 8'h28 ||
	       cpReq[11:4] == 8'h2C,
	       IF_cpReq_363_BITS_11_TO_4_366_EQ_0x0_445_THEN__ETC___d6178 } ;
  assign adminResp1F$ENQ = WILL_FIRE_RL_cpDispatch_F_T_T_T ;
  assign adminResp1F$DEQ =
	     WILL_FIRE_RL_readAdminResponseCollect && adminResp1F$EMPTY_N ;
  assign adminResp1F$CLR = 1'b0 ;

  // submodule adminResp2F
  always@(WILL_FIRE_RL_cpDispatch_F_T_T_F_T_T or
	  MUX_adminResp2F$enq_1__VAL_1 or
	  WILL_FIRE_RL_cpDispatch_F_T_T_F_T_F_T or
	  MUX_adminResp2F$enq_1__VAL_2 or
	  WILL_FIRE_RL_cpDispatch_F_T_T_F_T_F_F or
	  MUX_adminResp2F$enq_1__VAL_3)
  begin
    case (1'b1) // synopsys parallel_case
      WILL_FIRE_RL_cpDispatch_F_T_T_F_T_T:
	  adminResp2F$D_IN = MUX_adminResp2F$enq_1__VAL_1;
      WILL_FIRE_RL_cpDispatch_F_T_T_F_T_F_T:
	  adminResp2F$D_IN = MUX_adminResp2F$enq_1__VAL_2;
      WILL_FIRE_RL_cpDispatch_F_T_T_F_T_F_F:
	  adminResp2F$D_IN = MUX_adminResp2F$enq_1__VAL_3;
      default: adminResp2F$D_IN = 33'h0AAAAAAAA /* unspecified value */ ;
    endcase
  end
  assign adminResp2F$ENQ =
	     WILL_FIRE_RL_cpDispatch_F_T_T_F_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_T_T_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_T_T_F_T_F_F ;
  assign adminResp2F$DEQ =
	     WILL_FIRE_RL_readAdminResponseCollect && !adminResp1F$EMPTY_N &&
	     adminResp2F$EMPTY_N ;
  assign adminResp2F$CLR = 1'b0 ;

  // submodule adminResp3F
  assign adminResp3F$D_IN =
	     { cpReq[11:4] == 8'hC0 || cpReq[11:4] == 8'hC4 ||
	       cpReq[11:4] == 8'hC8 ||
	       cpReq[11:4] == 8'hCC ||
	       cpReq[11:4] == 8'hD0 ||
	       cpReq[11:4] == 8'hD4 ||
	       cpReq[11:4] == 8'hD8 ||
	       cpReq[11:4] == 8'hDC ||
	       cpReq[11:4] == 8'hE0 ||
	       cpReq[11:4] == 8'hE4 ||
	       cpReq[11:4] == 8'hE8 ||
	       cpReq[11:4] == 8'hEC ||
	       cpReq[11:4] == 8'hF0 ||
	       cpReq[11:4] == 8'hF4 ||
	       cpReq[11:4] == 8'hF8 ||
	       cpReq[11:4] == 8'hFC,
	       CASE_cpReq_BITS_9_TO_6_uuid_arg_BITS_31_TO_0_0_ETC__q3 } ;
  assign adminResp3F$ENQ = WILL_FIRE_RL_cpDispatch_F_T_T_F_F ;
  assign adminResp3F$DEQ =
	     WILL_FIRE_RL_readAdminResponseCollect && !adminResp1F$EMPTY_N &&
	     !adminResp2F$EMPTY_N &&
	     adminResp3F$EMPTY_N ;
  assign adminResp3F$CLR = 1'b0 ;

  // submodule adminResp4F
`ifdef not
  assign adminResp4F$D_IN = { 1'd1, rom_serverAdapter_outData_outData$wget } ;
  assign adminResp4F$ENQ = rom_serverAdapter_outData_deqCalled$whas ;
`else
  assign adminResp4F$D_IN = { 1'd1, 32'd0 } ;
  assign adminResp4F$ENQ = 1'b0 ;
`endif
  assign adminResp4F$DEQ =
	     WILL_FIRE_RL_readAdminResponseCollect && !adminResp1F$EMPTY_N &&
	     !adminResp2F$EMPTY_N &&
	     !adminResp3F$EMPTY_N &&
	     adminResp4F$EMPTY_N ;
  assign adminResp4F$CLR = 1'b0 ;
	      
  // submodule adminRespF
  assign adminRespF$D_IN =
	     adminResp1F$EMPTY_N ?
	       adminResp1F$D_OUT :
	       IF_adminResp2F_notEmpty__304_THEN_adminResp2F__ETC___d2342 ;
  assign adminRespF$ENQ =
	     WILL_FIRE_RL_readAdminResponseCollect &&
	     (adminResp1F$EMPTY_N || adminResp2F$EMPTY_N ||
	      adminResp3F$EMPTY_N ||
	      adminResp4F$EMPTY_N) ;
  assign adminRespF$DEQ = WILL_FIRE_RL_responseAdminRd ;
  assign adminRespF$CLR = 1'b0 ;

  // submodule cpReqF
  assign cpReqF$D_IN = server_request_put ;
  assign cpReqF$ENQ = EN_server_request_put ;
  assign cpReqF$DEQ = WILL_FIRE_RL_reqRcv ;
  assign cpReqF$CLR = 1'b0 ;

  // submodule cpRespF
  assign cpRespF$D_IN =
	     WILL_FIRE_RL_responseAdminRd ?
	       MUX_cpRespF$enq_1__VAL_1 :
	       MUX_cpRespF$enq_1__VAL_2 ;
  assign cpRespF$ENQ =
	     WILL_FIRE_RL_responseAdminRd || WILL_FIRE_RL_completeWorkerRead ;
  assign cpRespF$DEQ = EN_server_response_get ;
  assign cpRespF$CLR = 1'b0 ;

`ifdef not
  // submodule dna_dna
  assign dna_dna$CLK = dna_cnt[0] ;
  assign dna_dna$DIN = 1'd0 ;
  assign dna_dna$READ = dna_rdReg ;
  assign dna_dna$SHIFT = dna_shftReg ;

  // submodule rom_memory
  assign rom_memory$ADDR = cpReq[15:6] ;
  assign rom_memory$DI = 32'd0 ;
  assign rom_memory$WE = 1'd0 ;
  assign rom_memory$EN =
	     WILL_FIRE_RL_rom_serverAdapter_stageReadResponseAlways ;

  // submodule rom_serverAdapter_outDataCore
  assign rom_serverAdapter_outDataCore$D_IN = rom_memory$DO ;
  assign rom_serverAdapter_outDataCore$ENQ =
	     WILL_FIRE_RL_rom_serverAdapter_outData_enqAndDeq ||
	     rom_serverAdapter_outDataCore$FULL_N &&
	     !rom_serverAdapter_outData_deqCalled$whas &&
	     rom_serverAdapter_outData_enqData$whas ;
  assign rom_serverAdapter_outDataCore$DEQ =
	     WILL_FIRE_RL_rom_serverAdapter_outData_enqAndDeq ||
	     rom_serverAdapter_outDataCore$EMPTY_N &&
	     rom_serverAdapter_outData_deqCalled$whas &&
	     !rom_serverAdapter_outData_enqData$whas ;
  assign rom_serverAdapter_outDataCore$CLR = 1'b0 ;

  // submodule timeServ_disableServo
  assign timeServ_disableServo$sD_IN = timeServ_rplTimeControl[4] ;
  assign timeServ_disableServo$sEN = timeServ_disableServo$sRDY ;

  // submodule timeServ_nowInCC
  assign timeServ_nowInCC$sD_IN =
	     { timeServ_refSecCount, timeServ_fracSeconds[47:16] } ;
  assign timeServ_nowInCC$sEN = timeServ_nowInCC$sRDY ;

  // submodule timeServ_ppsDisablePPS
  assign timeServ_ppsDisablePPS$sD_IN = timeServ_rplTimeControl[2] ;
  assign timeServ_ppsDisablePPS$sEN = timeServ_ppsDisablePPS$sRDY ;

  // submodule timeServ_ppsLostCC
  assign timeServ_ppsLostCC$sD_IN = timeServ_ppsLost ;
  assign timeServ_ppsLostCC$sEN = timeServ_ppsLostCC$sRDY ;

  // submodule timeServ_ppsOKCC
  assign timeServ_ppsOKCC$sD_IN = timeServ_ppsOK ;
  assign timeServ_ppsOKCC$sEN = timeServ_ppsOKCC$sRDY ;

  // submodule timeServ_ppsOutMode
  assign timeServ_ppsOutMode$sD_IN = timeServ_rplTimeControl[1:0] ;
  assign timeServ_ppsOutMode$sEN = timeServ_ppsOutMode$sRDY ;

  // submodule timeServ_refPerPPS
  assign timeServ_refPerPPS$sD_IN = timeServ_refFreeSpan ;
  assign timeServ_refPerPPS$sEN =
	     timeServ_refPerPPS$sRDY && timeServ_ppsExtSync_d2 &&
	     !timeServ_ppsExtSyncD ;

  // submodule timeServ_rollingPPSIn
  assign timeServ_rollingPPSIn$sD_IN = timeServ_ppsEdgeCount ;
  assign timeServ_rollingPPSIn$sEN = timeServ_rollingPPSIn$sRDY ;

  // submodule timeServ_setRefF
  assign timeServ_setRefF$sD_IN = { td, cpReq[59:28] } ;
  assign timeServ_setRefF$sENQ = WILL_FIRE_RL_cpDispatch_T_F_F_F_F_F_F_T ;
  assign timeServ_setRefF$dDEQ = timeServ_setRefF$dEMPTY_N ;
`endif

  // submodule wci_mReset
  assign wci_mReset$ASSERT_IN = !wci_wReset_n ;

  // submodule wci_mReset_1
  assign wci_mReset_1$ASSERT_IN = !wci_wReset_n_1 ;

  // submodule wci_mReset_10
  assign wci_mReset_10$ASSERT_IN = !wci_wReset_n_10 ;

  // submodule wci_mReset_11
  assign wci_mReset_11$ASSERT_IN = !wci_wReset_n_11 ;

  // submodule wci_mReset_12
  assign wci_mReset_12$ASSERT_IN = !wci_wReset_n_12 ;

  // submodule wci_mReset_13
  assign wci_mReset_13$ASSERT_IN = !wci_wReset_n_13 ;

  // submodule wci_mReset_14
  assign wci_mReset_14$ASSERT_IN = !wci_wReset_n_14 ;

  // submodule wci_mReset_2
  assign wci_mReset_2$ASSERT_IN = !wci_wReset_n_2 ;

  // submodule wci_mReset_3
  assign wci_mReset_3$ASSERT_IN = !wci_wReset_n_3 ;

  // submodule wci_mReset_4
  assign wci_mReset_4$ASSERT_IN = !wci_wReset_n_4 ;

  // submodule wci_mReset_5
  assign wci_mReset_5$ASSERT_IN = !wci_wReset_n_5 ;

  // submodule wci_mReset_6
  assign wci_mReset_6$ASSERT_IN = !wci_wReset_n_6 ;

  // submodule wci_mReset_7
  assign wci_mReset_7$ASSERT_IN = !wci_wReset_n_7 ;

  // submodule wci_mReset_8
  assign wci_mReset_8$ASSERT_IN = !wci_wReset_n_8 ;

  // submodule wci_mReset_9
  assign wci_mReset_9$ASSERT_IN = !wci_wReset_n_9 ;

  // submodule wci_respF
  always@(MUX_wci_busy$write_1__SEL_1 or
	  MUX_wci_respF$enq_1__VAL_1 or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_T_F_F_T or
	  MUX_wci_respF$enq_1__VAL_2 or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_T_F_F_F_T or
	  MUX_wci_respF$enq_1__VAL_3 or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_T_F_F_F_F_T or
	  MUX_wci_respF$enq_1__VAL_4 or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_T_F_F_F_F_F_T or
	  MUX_wci_respF$enq_1__VAL_5 or
	  MUX_wci_respF$enq_1__SEL_6 or
	  MUX_wci_respF$enq_1__SEL_7 or WILL_FIRE_RL_cpDispatch_F_F_T_T_F_T)
  begin
    case (1'b1) // synopsys parallel_case
      MUX_wci_busy$write_1__SEL_1:
	  wci_respF$D_IN = MUX_wci_respF$enq_1__VAL_1;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_T_F_F_T:
	  wci_respF$D_IN = MUX_wci_respF$enq_1__VAL_2;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_T_F_F_F_T:
	  wci_respF$D_IN = MUX_wci_respF$enq_1__VAL_3;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_T_F_F_F_F_T:
	  wci_respF$D_IN = MUX_wci_respF$enq_1__VAL_4;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_T_F_F_F_F_F_T:
	  wci_respF$D_IN = MUX_wci_respF$enq_1__VAL_5;
      MUX_wci_respF$enq_1__SEL_6: wci_respF$D_IN = 34'h100000000;
      MUX_wci_respF$enq_1__SEL_7: wci_respF$D_IN = 34'h1C0DE4204;
      WILL_FIRE_RL_cpDispatch_F_F_T_T_F_T: wci_respF$D_IN = 34'h3C0DE4202;
      default: wci_respF$D_IN = 34'h2AAAAAAAA /* unspecified value */ ;
    endcase
  end
  assign wci_respF$ENQ =
	     WILL_FIRE_RL_wci_wrkBusy &&
	     (!wci_respTimr_28_ULT_1_SL_wci_wTimeout_29_30___d5879 ||
	      wci_wciResponse$wget[33:32] != 2'd0) ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_T_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_T_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_T_F_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_T_F_F_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_T_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_T_F_F_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_T_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_T_F_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_T_F_T ;
  assign wci_respF$DEQ = MUX_wrkAct$write_1__SEL_3 && wrkAct == 4'd0 ;
  assign wci_respF$CLR = 1'b0 ;

  // submodule wci_respF_1
  always@(MUX_wci_busy_1$write_1__SEL_1 or
	  MUX_wci_respF_1$enq_1__VAL_1 or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_F_F_T or
	  MUX_wci_respF_1$enq_1__VAL_2 or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_F_F_F_T or
	  MUX_wci_respF_1$enq_1__VAL_3 or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_F_F_F_F_T or
	  MUX_wci_respF_1$enq_1__VAL_4 or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_F_F_F_F_F_T or
	  MUX_wci_respF_1$enq_1__VAL_5 or
	  MUX_wci_respF_1$enq_1__SEL_6 or
	  MUX_wci_respF_1$enq_1__SEL_7 or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_T_F_T)
  begin
    case (1'b1) // synopsys parallel_case
      MUX_wci_busy_1$write_1__SEL_1:
	  wci_respF_1$D_IN = MUX_wci_respF_1$enq_1__VAL_1;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_F_F_T:
	  wci_respF_1$D_IN = MUX_wci_respF_1$enq_1__VAL_2;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_F_F_F_T:
	  wci_respF_1$D_IN = MUX_wci_respF_1$enq_1__VAL_3;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_F_F_F_F_T:
	  wci_respF_1$D_IN = MUX_wci_respF_1$enq_1__VAL_4;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_F_F_F_F_F_T:
	  wci_respF_1$D_IN = MUX_wci_respF_1$enq_1__VAL_5;
      MUX_wci_respF_1$enq_1__SEL_6: wci_respF_1$D_IN = 34'h100000000;
      MUX_wci_respF_1$enq_1__SEL_7: wci_respF_1$D_IN = 34'h1C0DE4204;
      WILL_FIRE_RL_cpDispatch_F_F_T_F_T_F_T: wci_respF_1$D_IN = 34'h3C0DE4202;
      default: wci_respF_1$D_IN = 34'h2AAAAAAAA /* unspecified value */ ;
    endcase
  end
  assign wci_respF_1$ENQ =
	     WILL_FIRE_RL_wci_wrkBusy_1 &&
	     (!wci_respTimr_1_68_ULT_1_SL_wci_wTimeout_1_69_70___d5880 ||
	      wci_wciResponse_1$wget[33:32] != 2'd0) ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_F_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_F_F_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_T_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_T_F_F_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_T_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_F_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_T_F_T ;
  assign wci_respF_1$DEQ = MUX_wrkAct$write_1__SEL_3 && wrkAct == 4'd1 ;
  assign wci_respF_1$CLR = 1'b0 ;

  // submodule wci_respF_10
  always@(MUX_wci_busy_10$write_1__SEL_1 or
	  MUX_wci_respF_10$enq_1__VAL_1 or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T or
	  MUX_wci_respF_10$enq_1__VAL_2 or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T or
	  MUX_wci_respF_10$enq_1__VAL_3 or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T or
	  MUX_wci_respF_10$enq_1__VAL_4 or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T or
	  MUX_wci_respF_10$enq_1__VAL_5 or
	  MUX_wci_respF_10$enq_1__SEL_6 or
	  MUX_wci_respF_10$enq_1__SEL_7 or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_T)
  begin
    case (1'b1) // synopsys parallel_case
      MUX_wci_busy_10$write_1__SEL_1:
	  wci_respF_10$D_IN = MUX_wci_respF_10$enq_1__VAL_1;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T:
	  wci_respF_10$D_IN = MUX_wci_respF_10$enq_1__VAL_2;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T:
	  wci_respF_10$D_IN = MUX_wci_respF_10$enq_1__VAL_3;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T:
	  wci_respF_10$D_IN = MUX_wci_respF_10$enq_1__VAL_4;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T:
	  wci_respF_10$D_IN = MUX_wci_respF_10$enq_1__VAL_5;
      MUX_wci_respF_10$enq_1__SEL_6: wci_respF_10$D_IN = 34'h100000000;
      MUX_wci_respF_10$enq_1__SEL_7: wci_respF_10$D_IN = 34'h1C0DE4204;
      WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_T:
	  wci_respF_10$D_IN = 34'h3C0DE4202;
      default: wci_respF_10$D_IN = 34'h2AAAAAAAA /* unspecified value */ ;
    endcase
  end
  assign wci_respF_10$ENQ =
	     WILL_FIRE_RL_wci_wrkBusy_10 &&
	     (!wci_respTimr_10_628_ULT_1_SL_wci_wTimeout_10_6_ETC___d5889 ||
	      wci_wciResponse_10$wget[33:32] != 2'd0) ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_T ;
  assign wci_respF_10$DEQ = MUX_wrkAct$write_1__SEL_3 && wrkAct == 4'd10 ;
  assign wci_respF_10$CLR = 1'b0 ;

  // submodule wci_respF_11
  always@(MUX_wci_busy_11$write_1__SEL_1 or
	  MUX_wci_respF_11$enq_1__VAL_1 or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T or
	  MUX_wci_respF_11$enq_1__VAL_2 or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T or
	  MUX_wci_respF_11$enq_1__VAL_3 or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T or
	  MUX_wci_respF_11$enq_1__VAL_4 or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T or
	  MUX_wci_respF_11$enq_1__VAL_5 or
	  MUX_wci_respF_11$enq_1__SEL_6 or
	  MUX_wci_respF_11$enq_1__SEL_7 or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_T)
  begin
    case (1'b1) // synopsys parallel_case
      MUX_wci_busy_11$write_1__SEL_1:
	  wci_respF_11$D_IN = MUX_wci_respF_11$enq_1__VAL_1;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T:
	  wci_respF_11$D_IN = MUX_wci_respF_11$enq_1__VAL_2;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T:
	  wci_respF_11$D_IN = MUX_wci_respF_11$enq_1__VAL_3;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T:
	  wci_respF_11$D_IN = MUX_wci_respF_11$enq_1__VAL_4;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T:
	  wci_respF_11$D_IN = MUX_wci_respF_11$enq_1__VAL_5;
      MUX_wci_respF_11$enq_1__SEL_6: wci_respF_11$D_IN = 34'h100000000;
      MUX_wci_respF_11$enq_1__SEL_7: wci_respF_11$D_IN = 34'h1C0DE4204;
      WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_T:
	  wci_respF_11$D_IN = 34'h3C0DE4202;
      default: wci_respF_11$D_IN = 34'h2AAAAAAAA /* unspecified value */ ;
    endcase
  end
  assign wci_respF_11$ENQ =
	     WILL_FIRE_RL_wci_wrkBusy_11 &&
	     (!wci_respTimr_11_768_ULT_1_SL_wci_wTimeout_11_7_ETC___d5890 ||
	      wci_wciResponse_11$wget[33:32] != 2'd0) ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_T ;
  assign wci_respF_11$DEQ = MUX_wrkAct$write_1__SEL_3 && wrkAct == 4'd11 ;
  assign wci_respF_11$CLR = 1'b0 ;

  // submodule wci_respF_12
  always@(MUX_wci_busy_12$write_1__SEL_1 or
	  MUX_wci_respF_12$enq_1__VAL_1 or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T or
	  MUX_wci_respF_12$enq_1__VAL_2 or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T or
	  MUX_wci_respF_12$enq_1__VAL_3 or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T or
	  MUX_wci_respF_12$enq_1__VAL_4 or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T or
	  MUX_wci_respF_12$enq_1__VAL_5 or
	  MUX_wci_respF_12$enq_1__SEL_6 or
	  MUX_wci_respF_12$enq_1__SEL_7 or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T)
  begin
    case (1'b1) // synopsys parallel_case
      MUX_wci_busy_12$write_1__SEL_1:
	  wci_respF_12$D_IN = MUX_wci_respF_12$enq_1__VAL_1;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T:
	  wci_respF_12$D_IN = MUX_wci_respF_12$enq_1__VAL_2;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T:
	  wci_respF_12$D_IN = MUX_wci_respF_12$enq_1__VAL_3;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T:
	  wci_respF_12$D_IN = MUX_wci_respF_12$enq_1__VAL_4;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T:
	  wci_respF_12$D_IN = MUX_wci_respF_12$enq_1__VAL_5;
      MUX_wci_respF_12$enq_1__SEL_6: wci_respF_12$D_IN = 34'h100000000;
      MUX_wci_respF_12$enq_1__SEL_7: wci_respF_12$D_IN = 34'h1C0DE4204;
      WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T:
	  wci_respF_12$D_IN = 34'h3C0DE4202;
      default: wci_respF_12$D_IN = 34'h2AAAAAAAA /* unspecified value */ ;
    endcase
  end
  assign wci_respF_12$ENQ =
	     WILL_FIRE_RL_wci_wrkBusy_12 &&
	     (!wci_respTimr_12_908_ULT_1_SL_wci_wTimeout_12_9_ETC___d5891 ||
	      wci_wciResponse_12$wget[33:32] != 2'd0) ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T ;
  assign wci_respF_12$DEQ = MUX_wrkAct$write_1__SEL_3 && wrkAct == 4'd12 ;
  assign wci_respF_12$CLR = 1'b0 ;

  // submodule wci_respF_13
  always@(MUX_wci_busy_13$write_1__SEL_1 or
	  MUX_wci_respF_13$enq_1__VAL_1 or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T or
	  MUX_wci_respF_13$enq_1__VAL_2 or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T or
	  MUX_wci_respF_13$enq_1__VAL_3 or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T or
	  MUX_wci_respF_13$enq_1__VAL_4 or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T or
	  MUX_wci_respF_13$enq_1__VAL_5 or
	  MUX_wci_respF_13$enq_1__SEL_6 or
	  MUX_wci_respF_13$enq_1__SEL_7 or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T)
  begin
    case (1'b1) // synopsys parallel_case
      MUX_wci_busy_13$write_1__SEL_1:
	  wci_respF_13$D_IN = MUX_wci_respF_13$enq_1__VAL_1;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T:
	  wci_respF_13$D_IN = MUX_wci_respF_13$enq_1__VAL_2;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T:
	  wci_respF_13$D_IN = MUX_wci_respF_13$enq_1__VAL_3;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T:
	  wci_respF_13$D_IN = MUX_wci_respF_13$enq_1__VAL_4;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T:
	  wci_respF_13$D_IN = MUX_wci_respF_13$enq_1__VAL_5;
      MUX_wci_respF_13$enq_1__SEL_6: wci_respF_13$D_IN = 34'h100000000;
      MUX_wci_respF_13$enq_1__SEL_7: wci_respF_13$D_IN = 34'h1C0DE4204;
      WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T:
	  wci_respF_13$D_IN = 34'h3C0DE4202;
      default: wci_respF_13$D_IN = 34'h2AAAAAAAA /* unspecified value */ ;
    endcase
  end
  assign wci_respF_13$ENQ =
	     WILL_FIRE_RL_wci_wrkBusy_13 &&
	     (!wci_respTimr_13_048_ULT_1_SL_wci_wTimeout_13_0_ETC___d5892 ||
	      wci_wciResponse_13$wget[33:32] != 2'd0) ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T ;
  assign wci_respF_13$DEQ = MUX_wrkAct$write_1__SEL_3 && wrkAct == 4'd13 ;
  assign wci_respF_13$CLR = 1'b0 ;

  // submodule wci_respF_14
  always@(MUX_wci_busy_14$write_1__SEL_1 or
	  MUX_wci_respF_14$enq_1__VAL_1 or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T or
	  MUX_wci_respF_14$enq_1__VAL_2 or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T or
	  MUX_wci_respF_14$enq_1__VAL_3 or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T or
	  MUX_wci_respF_14$enq_1__VAL_4 or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T or
	  MUX_wci_respF_14$enq_1__VAL_5 or
	  MUX_wci_respF_14$enq_1__SEL_6 or
	  MUX_wci_respF_14$enq_1__SEL_7 or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T)
  begin
    case (1'b1) // synopsys parallel_case
      MUX_wci_busy_14$write_1__SEL_1:
	  wci_respF_14$D_IN = MUX_wci_respF_14$enq_1__VAL_1;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T:
	  wci_respF_14$D_IN = MUX_wci_respF_14$enq_1__VAL_2;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T:
	  wci_respF_14$D_IN = MUX_wci_respF_14$enq_1__VAL_3;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T:
	  wci_respF_14$D_IN = MUX_wci_respF_14$enq_1__VAL_4;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T:
	  wci_respF_14$D_IN = MUX_wci_respF_14$enq_1__VAL_5;
      MUX_wci_respF_14$enq_1__SEL_6: wci_respF_14$D_IN = 34'h100000000;
      MUX_wci_respF_14$enq_1__SEL_7: wci_respF_14$D_IN = 34'h1C0DE4204;
      WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T:
	  wci_respF_14$D_IN = 34'h3C0DE4202;
      default: wci_respF_14$D_IN = 34'h2AAAAAAAA /* unspecified value */ ;
    endcase
  end
  assign wci_respF_14$ENQ =
	     WILL_FIRE_RL_wci_wrkBusy_14 &&
	     (!wci_respTimr_14_188_ULT_1_SL_wci_wTimeout_14_1_ETC___d5893 ||
	      wci_wciResponse_14$wget[33:32] != 2'd0) ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T ;
  assign wci_respF_14$DEQ = MUX_wrkAct$write_1__SEL_3 && wrkAct == 4'd14 ;
  assign wci_respF_14$CLR = 1'b0 ;

  // submodule wci_respF_2
  always@(MUX_wci_busy_2$write_1__SEL_1 or
	  MUX_wci_respF_2$enq_1__VAL_1 or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_F_F_T or
	  MUX_wci_respF_2$enq_1__VAL_2 or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_F_F_F_T or
	  MUX_wci_respF_2$enq_1__VAL_3 or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_F_F_F_F_T or
	  MUX_wci_respF_2$enq_1__VAL_4 or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_F_F_F_F_F_T or
	  MUX_wci_respF_2$enq_1__VAL_5 or
	  MUX_wci_respF_2$enq_1__SEL_6 or
	  MUX_wci_respF_2$enq_1__SEL_7 or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_F_T)
  begin
    case (1'b1) // synopsys parallel_case
      MUX_wci_busy_2$write_1__SEL_1:
	  wci_respF_2$D_IN = MUX_wci_respF_2$enq_1__VAL_1;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_F_F_T:
	  wci_respF_2$D_IN = MUX_wci_respF_2$enq_1__VAL_2;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_F_F_F_T:
	  wci_respF_2$D_IN = MUX_wci_respF_2$enq_1__VAL_3;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_F_F_F_F_T:
	  wci_respF_2$D_IN = MUX_wci_respF_2$enq_1__VAL_4;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_F_F_F_F_F_T:
	  wci_respF_2$D_IN = MUX_wci_respF_2$enq_1__VAL_5;
      MUX_wci_respF_2$enq_1__SEL_6: wci_respF_2$D_IN = 34'h100000000;
      MUX_wci_respF_2$enq_1__SEL_7: wci_respF_2$D_IN = 34'h1C0DE4204;
      WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_F_T:
	  wci_respF_2$D_IN = 34'h3C0DE4202;
      default: wci_respF_2$D_IN = 34'h2AAAAAAAA /* unspecified value */ ;
    endcase
  end
  assign wci_respF_2$ENQ =
	     WILL_FIRE_RL_wci_wrkBusy_2 &&
	     (!wci_respTimr_2_08_ULT_1_SL_wci_wTimeout_2_09_10___d5881 ||
	      wci_wciResponse_2$wget[33:32] != 2'd0) ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_F_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_F_F_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_F_F_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_F_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_F_T ;
  assign wci_respF_2$DEQ = MUX_wrkAct$write_1__SEL_3 && wrkAct == 4'd2 ;
  assign wci_respF_2$CLR = 1'b0 ;

  // submodule wci_respF_3
  always@(MUX_wci_busy_3$write_1__SEL_1 or
	  MUX_wci_respF_3$enq_1__VAL_1 or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_F_F_T or
	  MUX_wci_respF_3$enq_1__VAL_2 or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_F_F_F_T or
	  MUX_wci_respF_3$enq_1__VAL_3 or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_F_F_F_F_T or
	  MUX_wci_respF_3$enq_1__VAL_4 or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_F_F_F_F_F_T or
	  MUX_wci_respF_3$enq_1__VAL_5 or
	  MUX_wci_respF_3$enq_1__SEL_6 or
	  MUX_wci_respF_3$enq_1__SEL_7 or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_F_T)
  begin
    case (1'b1) // synopsys parallel_case
      MUX_wci_busy_3$write_1__SEL_1:
	  wci_respF_3$D_IN = MUX_wci_respF_3$enq_1__VAL_1;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_F_F_T:
	  wci_respF_3$D_IN = MUX_wci_respF_3$enq_1__VAL_2;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_F_F_F_T:
	  wci_respF_3$D_IN = MUX_wci_respF_3$enq_1__VAL_3;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_F_F_F_F_T:
	  wci_respF_3$D_IN = MUX_wci_respF_3$enq_1__VAL_4;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_F_F_F_F_F_T:
	  wci_respF_3$D_IN = MUX_wci_respF_3$enq_1__VAL_5;
      MUX_wci_respF_3$enq_1__SEL_6: wci_respF_3$D_IN = 34'h100000000;
      MUX_wci_respF_3$enq_1__SEL_7: wci_respF_3$D_IN = 34'h1C0DE4204;
      WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_F_T:
	  wci_respF_3$D_IN = 34'h3C0DE4202;
      default: wci_respF_3$D_IN = 34'h2AAAAAAAA /* unspecified value */ ;
    endcase
  end
  assign wci_respF_3$ENQ =
	     WILL_FIRE_RL_wci_wrkBusy_3 &&
	     (!wci_respTimr_3_48_ULT_1_SL_wci_wTimeout_3_49_50___d5882 ||
	      wci_wciResponse_3$wget[33:32] != 2'd0) ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_F_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_F_F_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_F_F_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_F_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_F_T ;
  assign wci_respF_3$DEQ = MUX_wrkAct$write_1__SEL_3 && wrkAct == 4'd3 ;
  assign wci_respF_3$CLR = 1'b0 ;

  // submodule wci_respF_4
  always@(MUX_wci_busy_4$write_1__SEL_1 or
	  MUX_wci_respF_4$enq_1__VAL_1 or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_F_F_T or
	  MUX_wci_respF_4$enq_1__VAL_2 or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_F_F_F_T or
	  MUX_wci_respF_4$enq_1__VAL_3 or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_F_F_F_F_T or
	  MUX_wci_respF_4$enq_1__VAL_4 or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T or
	  MUX_wci_respF_4$enq_1__VAL_5 or
	  MUX_wci_respF_4$enq_1__SEL_6 or
	  MUX_wci_respF_4$enq_1__SEL_7 or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_F_T)
  begin
    case (1'b1) // synopsys parallel_case
      MUX_wci_busy_4$write_1__SEL_1:
	  wci_respF_4$D_IN = MUX_wci_respF_4$enq_1__VAL_1;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_F_F_T:
	  wci_respF_4$D_IN = MUX_wci_respF_4$enq_1__VAL_2;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_F_F_F_T:
	  wci_respF_4$D_IN = MUX_wci_respF_4$enq_1__VAL_3;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_F_F_F_F_T:
	  wci_respF_4$D_IN = MUX_wci_respF_4$enq_1__VAL_4;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T:
	  wci_respF_4$D_IN = MUX_wci_respF_4$enq_1__VAL_5;
      MUX_wci_respF_4$enq_1__SEL_6: wci_respF_4$D_IN = 34'h100000000;
      MUX_wci_respF_4$enq_1__SEL_7: wci_respF_4$D_IN = 34'h1C0DE4204;
      WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_F_T:
	  wci_respF_4$D_IN = 34'h3C0DE4202;
      default: wci_respF_4$D_IN = 34'h2AAAAAAAA /* unspecified value */ ;
    endcase
  end
  assign wci_respF_4$ENQ =
	     WILL_FIRE_RL_wci_wrkBusy_4 &&
	     (!wci_respTimr_4_88_ULT_1_SL_wci_wTimeout_4_89_90___d5883 ||
	      wci_wciResponse_4$wget[33:32] != 2'd0) ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_F_F_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_F_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_F_T ;
  assign wci_respF_4$DEQ = MUX_wrkAct$write_1__SEL_3 && wrkAct == 4'd4 ;
  assign wci_respF_4$CLR = 1'b0 ;

  // submodule wci_respF_5
  always@(MUX_wci_busy_5$write_1__SEL_1 or
	  MUX_wci_respF_5$enq_1__VAL_1 or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_F_F_T or
	  MUX_wci_respF_5$enq_1__VAL_2 or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_F_F_F_T or
	  MUX_wci_respF_5$enq_1__VAL_3 or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T or
	  MUX_wci_respF_5$enq_1__VAL_4 or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T or
	  MUX_wci_respF_5$enq_1__VAL_5 or
	  MUX_wci_respF_5$enq_1__SEL_6 or
	  MUX_wci_respF_5$enq_1__SEL_7 or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_T)
  begin
    case (1'b1) // synopsys parallel_case
      MUX_wci_busy_5$write_1__SEL_1:
	  wci_respF_5$D_IN = MUX_wci_respF_5$enq_1__VAL_1;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_F_F_T:
	  wci_respF_5$D_IN = MUX_wci_respF_5$enq_1__VAL_2;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_F_F_F_T:
	  wci_respF_5$D_IN = MUX_wci_respF_5$enq_1__VAL_3;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T:
	  wci_respF_5$D_IN = MUX_wci_respF_5$enq_1__VAL_4;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T:
	  wci_respF_5$D_IN = MUX_wci_respF_5$enq_1__VAL_5;
      MUX_wci_respF_5$enq_1__SEL_6: wci_respF_5$D_IN = 34'h100000000;
      MUX_wci_respF_5$enq_1__SEL_7: wci_respF_5$D_IN = 34'h1C0DE4204;
      WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_T:
	  wci_respF_5$D_IN = 34'h3C0DE4202;
      default: wci_respF_5$D_IN = 34'h2AAAAAAAA /* unspecified value */ ;
    endcase
  end
  assign wci_respF_5$ENQ =
	     WILL_FIRE_RL_wci_wrkBusy_5 &&
	     (!wci_respTimr_5_28_ULT_1_SL_wci_wTimeout_5_29_30___d5884 ||
	      wci_wciResponse_5$wget[33:32] != 2'd0) ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_F_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_F_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_T ;
  assign wci_respF_5$DEQ = MUX_wrkAct$write_1__SEL_3 && wrkAct == 4'd5 ;
  assign wci_respF_5$CLR = 1'b0 ;

  // submodule wci_respF_6
  always@(MUX_wci_busy_6$write_1__SEL_1 or
	  MUX_wci_respF_6$enq_1__VAL_1 or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_F_F_T or
	  MUX_wci_respF_6$enq_1__VAL_2 or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T or
	  MUX_wci_respF_6$enq_1__VAL_3 or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T or
	  MUX_wci_respF_6$enq_1__VAL_4 or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T or
	  MUX_wci_respF_6$enq_1__VAL_5 or
	  MUX_wci_respF_6$enq_1__SEL_6 or
	  MUX_wci_respF_6$enq_1__SEL_7 or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_T)
  begin
    case (1'b1) // synopsys parallel_case
      MUX_wci_busy_6$write_1__SEL_1:
	  wci_respF_6$D_IN = MUX_wci_respF_6$enq_1__VAL_1;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_F_F_T:
	  wci_respF_6$D_IN = MUX_wci_respF_6$enq_1__VAL_2;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T:
	  wci_respF_6$D_IN = MUX_wci_respF_6$enq_1__VAL_3;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T:
	  wci_respF_6$D_IN = MUX_wci_respF_6$enq_1__VAL_4;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T:
	  wci_respF_6$D_IN = MUX_wci_respF_6$enq_1__VAL_5;
      MUX_wci_respF_6$enq_1__SEL_6: wci_respF_6$D_IN = 34'h100000000;
      MUX_wci_respF_6$enq_1__SEL_7: wci_respF_6$D_IN = 34'h1C0DE4204;
      WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_T:
	  wci_respF_6$D_IN = 34'h3C0DE4202;
      default: wci_respF_6$D_IN = 34'h2AAAAAAAA /* unspecified value */ ;
    endcase
  end
  assign wci_respF_6$ENQ =
	     WILL_FIRE_RL_wci_wrkBusy_6 &&
	     (!wci_respTimr_6_068_ULT_1_SL_wci_wTimeout_6_069_ETC___d5885 ||
	      wci_wciResponse_6$wget[33:32] != 2'd0) ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_F_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_F_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_T ;
  assign wci_respF_6$DEQ = MUX_wrkAct$write_1__SEL_3 && wrkAct == 4'd6 ;
  assign wci_respF_6$CLR = 1'b0 ;

  // submodule wci_respF_7
  always@(MUX_wci_busy_7$write_1__SEL_1 or
	  MUX_wci_respF_7$enq_1__VAL_1 or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T or
	  MUX_wci_respF_7$enq_1__VAL_2 or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T or
	  MUX_wci_respF_7$enq_1__VAL_3 or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T or
	  MUX_wci_respF_7$enq_1__VAL_4 or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T or
	  MUX_wci_respF_7$enq_1__VAL_5 or
	  MUX_wci_respF_7$enq_1__SEL_6 or
	  MUX_wci_respF_7$enq_1__SEL_7 or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_T)
  begin
    case (1'b1) // synopsys parallel_case
      MUX_wci_busy_7$write_1__SEL_1:
	  wci_respF_7$D_IN = MUX_wci_respF_7$enq_1__VAL_1;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T:
	  wci_respF_7$D_IN = MUX_wci_respF_7$enq_1__VAL_2;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T:
	  wci_respF_7$D_IN = MUX_wci_respF_7$enq_1__VAL_3;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T:
	  wci_respF_7$D_IN = MUX_wci_respF_7$enq_1__VAL_4;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T:
	  wci_respF_7$D_IN = MUX_wci_respF_7$enq_1__VAL_5;
      MUX_wci_respF_7$enq_1__SEL_6: wci_respF_7$D_IN = 34'h100000000;
      MUX_wci_respF_7$enq_1__SEL_7: wci_respF_7$D_IN = 34'h1C0DE4204;
      WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_T:
	  wci_respF_7$D_IN = 34'h3C0DE4202;
      default: wci_respF_7$D_IN = 34'h2AAAAAAAA /* unspecified value */ ;
    endcase
  end
  assign wci_respF_7$ENQ =
	     WILL_FIRE_RL_wci_wrkBusy_7 &&
	     (!wci_respTimr_7_208_ULT_1_SL_wci_wTimeout_7_209_ETC___d5886 ||
	      wci_wciResponse_7$wget[33:32] != 2'd0) ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_F_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_T ;
  assign wci_respF_7$DEQ = MUX_wrkAct$write_1__SEL_3 && wrkAct == 4'd7 ;
  assign wci_respF_7$CLR = 1'b0 ;

  // submodule wci_respF_8
  always@(MUX_wci_busy_8$write_1__SEL_1 or
	  MUX_wci_respF_8$enq_1__VAL_1 or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T or
	  MUX_wci_respF_8$enq_1__VAL_2 or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T or
	  MUX_wci_respF_8$enq_1__VAL_3 or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T or
	  MUX_wci_respF_8$enq_1__VAL_4 or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T or
	  MUX_wci_respF_8$enq_1__VAL_5 or
	  MUX_wci_respF_8$enq_1__SEL_6 or
	  MUX_wci_respF_8$enq_1__SEL_7 or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_T)
  begin
    case (1'b1) // synopsys parallel_case
      MUX_wci_busy_8$write_1__SEL_1:
	  wci_respF_8$D_IN = MUX_wci_respF_8$enq_1__VAL_1;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T:
	  wci_respF_8$D_IN = MUX_wci_respF_8$enq_1__VAL_2;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T:
	  wci_respF_8$D_IN = MUX_wci_respF_8$enq_1__VAL_3;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T:
	  wci_respF_8$D_IN = MUX_wci_respF_8$enq_1__VAL_4;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T:
	  wci_respF_8$D_IN = MUX_wci_respF_8$enq_1__VAL_5;
      MUX_wci_respF_8$enq_1__SEL_6: wci_respF_8$D_IN = 34'h100000000;
      MUX_wci_respF_8$enq_1__SEL_7: wci_respF_8$D_IN = 34'h1C0DE4204;
      WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_T:
	  wci_respF_8$D_IN = 34'h3C0DE4202;
      default: wci_respF_8$D_IN = 34'h2AAAAAAAA /* unspecified value */ ;
    endcase
  end
  assign wci_respF_8$ENQ =
	     WILL_FIRE_RL_wci_wrkBusy_8 &&
	     (!wci_respTimr_8_348_ULT_1_SL_wci_wTimeout_8_349_ETC___d5887 ||
	      wci_wciResponse_8$wget[33:32] != 2'd0) ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_F_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_T ;
  assign wci_respF_8$DEQ = MUX_wrkAct$write_1__SEL_3 && wrkAct == 4'd8 ;
  assign wci_respF_8$CLR = 1'b0 ;

  // submodule wci_respF_9
  always@(MUX_wci_busy_9$write_1__SEL_1 or
	  MUX_wci_respF_9$enq_1__VAL_1 or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T or
	  MUX_wci_respF_9$enq_1__VAL_2 or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T or
	  MUX_wci_respF_9$enq_1__VAL_3 or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T or
	  MUX_wci_respF_9$enq_1__VAL_4 or
	  WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T or
	  MUX_wci_respF_9$enq_1__VAL_5 or
	  MUX_wci_respF_9$enq_1__SEL_6 or
	  MUX_wci_respF_9$enq_1__SEL_7 or
	  WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_T)
  begin
    case (1'b1) // synopsys parallel_case
      MUX_wci_busy_9$write_1__SEL_1:
	  wci_respF_9$D_IN = MUX_wci_respF_9$enq_1__VAL_1;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T:
	  wci_respF_9$D_IN = MUX_wci_respF_9$enq_1__VAL_2;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T:
	  wci_respF_9$D_IN = MUX_wci_respF_9$enq_1__VAL_3;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T:
	  wci_respF_9$D_IN = MUX_wci_respF_9$enq_1__VAL_4;
      WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T:
	  wci_respF_9$D_IN = MUX_wci_respF_9$enq_1__VAL_5;
      MUX_wci_respF_9$enq_1__SEL_6: wci_respF_9$D_IN = 34'h100000000;
      MUX_wci_respF_9$enq_1__SEL_7: wci_respF_9$D_IN = 34'h1C0DE4204;
      WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_T:
	  wci_respF_9$D_IN = 34'h3C0DE4202;
      default: wci_respF_9$D_IN = 34'h2AAAAAAAA /* unspecified value */ ;
    endcase
  end
  assign wci_respF_9$ENQ =
	     WILL_FIRE_RL_wci_wrkBusy_9 &&
	     (!wci_respTimr_9_488_ULT_1_SL_wci_wTimeout_9_489_ETC___d5888 ||
	      wci_wciResponse_9$wget[33:32] != 2'd0) ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_F_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_F_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_F_T_F_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_F_T_F_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_T_F ||
	     WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_T ;
  assign wci_respF_9$DEQ = MUX_wrkAct$write_1__SEL_3 && wrkAct == 4'd9 ;
  assign wci_respF_9$CLR = 1'b0 ;

  // remaining internal signals
  assign IF_adminResp2F_notEmpty__304_THEN_adminResp2F__ETC___d2342 =
	     adminResp2F$EMPTY_N ?
	       adminResp2F$D_OUT :
	       (adminResp3F$EMPTY_N ? adminResp3F$D_OUT : adminResp4F$D_OUT) ;
  assign IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d3932 =
	     _theResult_____1__h76814 == 4'd0 && cpReq[37:36] != 2'd2 &&
	     cpReq[9:6] == 4'h8 &&
	     !wci_busy &&
	     wci_respF$FULL_N &&
	     !dispatched ;
  assign IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d3941 =
	     _theResult_____1__h76814 == 4'd0 && cpReq[37:36] != 2'd2 &&
	     cpReq[9:6] == 4'h9 &&
	     !wci_busy &&
	     wci_respF$FULL_N &&
	     !dispatched ;
  assign IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d3951 =
	     _theResult_____1__h76814 == 4'd0 && cpReq[37:36] != 2'd2 &&
	     cpReq[9:6] == 4'hA &&
	     !wci_busy &&
	     wci_respF$FULL_N &&
	     !dispatched ;
  assign IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4010 =
	     _theResult_____1__h76814 == 4'd1 && cpReq[37:36] != 2'd2 &&
	     cpReq[9:6] == 4'h8 &&
	     !wci_busy_1 &&
	     wci_respF_1$FULL_N &&
	     !dispatched ;
  assign IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4019 =
	     _theResult_____1__h76814 == 4'd1 && cpReq[37:36] != 2'd2 &&
	     cpReq[9:6] == 4'h9 &&
	     !wci_busy_1 &&
	     wci_respF_1$FULL_N &&
	     !dispatched ;
  assign IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4029 =
	     _theResult_____1__h76814 == 4'd1 && cpReq[37:36] != 2'd2 &&
	     cpReq[9:6] == 4'hA &&
	     !wci_busy_1 &&
	     wci_respF_1$FULL_N &&
	     !dispatched ;
  assign IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4086 =
	     _theResult_____1__h76814 == 4'd2 && cpReq[37:36] != 2'd2 &&
	     cpReq[9:6] == 4'h8 &&
	     !wci_busy_2 &&
	     wci_respF_2$FULL_N &&
	     !dispatched ;
  assign IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4095 =
	     _theResult_____1__h76814 == 4'd2 && cpReq[37:36] != 2'd2 &&
	     cpReq[9:6] == 4'h9 &&
	     !wci_busy_2 &&
	     wci_respF_2$FULL_N &&
	     !dispatched ;
  assign IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4105 =
	     _theResult_____1__h76814 == 4'd2 && cpReq[37:36] != 2'd2 &&
	     cpReq[9:6] == 4'hA &&
	     !wci_busy_2 &&
	     wci_respF_2$FULL_N &&
	     !dispatched ;
  assign IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4162 =
	     _theResult_____1__h76814 == 4'd3 && cpReq[37:36] != 2'd2 &&
	     cpReq[9:6] == 4'h8 &&
	     !wci_busy_3 &&
	     wci_respF_3$FULL_N &&
	     !dispatched ;
  assign IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4171 =
	     _theResult_____1__h76814 == 4'd3 && cpReq[37:36] != 2'd2 &&
	     cpReq[9:6] == 4'h9 &&
	     !wci_busy_3 &&
	     wci_respF_3$FULL_N &&
	     !dispatched ;
  assign IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4181 =
	     _theResult_____1__h76814 == 4'd3 && cpReq[37:36] != 2'd2 &&
	     cpReq[9:6] == 4'hA &&
	     !wci_busy_3 &&
	     wci_respF_3$FULL_N &&
	     !dispatched ;
  assign IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4238 =
	     _theResult_____1__h76814 == 4'd4 && cpReq[37:36] != 2'd2 &&
	     cpReq[9:6] == 4'h8 &&
	     !wci_busy_4 &&
	     wci_respF_4$FULL_N &&
	     !dispatched ;
  assign IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4247 =
	     _theResult_____1__h76814 == 4'd4 && cpReq[37:36] != 2'd2 &&
	     cpReq[9:6] == 4'h9 &&
	     !wci_busy_4 &&
	     wci_respF_4$FULL_N &&
	     !dispatched ;
  assign IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4257 =
	     _theResult_____1__h76814 == 4'd4 && cpReq[37:36] != 2'd2 &&
	     cpReq[9:6] == 4'hA &&
	     !wci_busy_4 &&
	     wci_respF_4$FULL_N &&
	     !dispatched ;
  assign IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4314 =
	     _theResult_____1__h76814 == 4'd5 && cpReq[37:36] != 2'd2 &&
	     cpReq[9:6] == 4'h8 &&
	     !wci_busy_5 &&
	     wci_respF_5$FULL_N &&
	     !dispatched ;
  assign IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4323 =
	     _theResult_____1__h76814 == 4'd5 && cpReq[37:36] != 2'd2 &&
	     cpReq[9:6] == 4'h9 &&
	     !wci_busy_5 &&
	     wci_respF_5$FULL_N &&
	     !dispatched ;
  assign IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4333 =
	     _theResult_____1__h76814 == 4'd5 && cpReq[37:36] != 2'd2 &&
	     cpReq[9:6] == 4'hA &&
	     !wci_busy_5 &&
	     wci_respF_5$FULL_N &&
	     !dispatched ;
  assign IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4390 =
	     _theResult_____1__h76814 == 4'd6 && cpReq[37:36] != 2'd2 &&
	     cpReq[9:6] == 4'h8 &&
	     !wci_busy_6 &&
	     wci_respF_6$FULL_N &&
	     !dispatched ;
  assign IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4399 =
	     _theResult_____1__h76814 == 4'd6 && cpReq[37:36] != 2'd2 &&
	     cpReq[9:6] == 4'h9 &&
	     !wci_busy_6 &&
	     wci_respF_6$FULL_N &&
	     !dispatched ;
  assign IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4409 =
	     _theResult_____1__h76814 == 4'd6 && cpReq[37:36] != 2'd2 &&
	     cpReq[9:6] == 4'hA &&
	     !wci_busy_6 &&
	     wci_respF_6$FULL_N &&
	     !dispatched ;
  assign IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4466 =
	     _theResult_____1__h76814 == 4'd7 && cpReq[37:36] != 2'd2 &&
	     cpReq[9:6] == 4'h8 &&
	     !wci_busy_7 &&
	     wci_respF_7$FULL_N &&
	     !dispatched ;
  assign IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4475 =
	     _theResult_____1__h76814 == 4'd7 && cpReq[37:36] != 2'd2 &&
	     cpReq[9:6] == 4'h9 &&
	     !wci_busy_7 &&
	     wci_respF_7$FULL_N &&
	     !dispatched ;
  assign IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4485 =
	     _theResult_____1__h76814 == 4'd7 && cpReq[37:36] != 2'd2 &&
	     cpReq[9:6] == 4'hA &&
	     !wci_busy_7 &&
	     wci_respF_7$FULL_N &&
	     !dispatched ;
  assign IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4542 =
	     _theResult_____1__h76814 == 4'd8 && cpReq[37:36] != 2'd2 &&
	     cpReq[9:6] == 4'h8 &&
	     !wci_busy_8 &&
	     wci_respF_8$FULL_N &&
	     !dispatched ;
  assign IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4551 =
	     _theResult_____1__h76814 == 4'd8 && cpReq[37:36] != 2'd2 &&
	     cpReq[9:6] == 4'h9 &&
	     !wci_busy_8 &&
	     wci_respF_8$FULL_N &&
	     !dispatched ;
  assign IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4561 =
	     _theResult_____1__h76814 == 4'd8 && cpReq[37:36] != 2'd2 &&
	     cpReq[9:6] == 4'hA &&
	     !wci_busy_8 &&
	     wci_respF_8$FULL_N &&
	     !dispatched ;
  assign IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4618 =
	     _theResult_____1__h76814 == 4'd9 && cpReq[37:36] != 2'd2 &&
	     cpReq[9:6] == 4'h8 &&
	     !wci_busy_9 &&
	     wci_respF_9$FULL_N &&
	     !dispatched ;
  assign IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4627 =
	     _theResult_____1__h76814 == 4'd9 && cpReq[37:36] != 2'd2 &&
	     cpReq[9:6] == 4'h9 &&
	     !wci_busy_9 &&
	     wci_respF_9$FULL_N &&
	     !dispatched ;
  assign IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4637 =
	     _theResult_____1__h76814 == 4'd9 && cpReq[37:36] != 2'd2 &&
	     cpReq[9:6] == 4'hA &&
	     !wci_busy_9 &&
	     wci_respF_9$FULL_N &&
	     !dispatched ;
  assign IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4694 =
	     _theResult_____1__h76814 == 4'd10 && cpReq[37:36] != 2'd2 &&
	     cpReq[9:6] == 4'h8 &&
	     !wci_busy_10 &&
	     wci_respF_10$FULL_N &&
	     !dispatched ;
  assign IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4703 =
	     _theResult_____1__h76814 == 4'd10 && cpReq[37:36] != 2'd2 &&
	     cpReq[9:6] == 4'h9 &&
	     !wci_busy_10 &&
	     wci_respF_10$FULL_N &&
	     !dispatched ;
  assign IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4713 =
	     _theResult_____1__h76814 == 4'd10 && cpReq[37:36] != 2'd2 &&
	     cpReq[9:6] == 4'hA &&
	     !wci_busy_10 &&
	     wci_respF_10$FULL_N &&
	     !dispatched ;
  assign IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4770 =
	     _theResult_____1__h76814 == 4'd11 && cpReq[37:36] != 2'd2 &&
	     cpReq[9:6] == 4'h8 &&
	     !wci_busy_11 &&
	     wci_respF_11$FULL_N &&
	     !dispatched ;
  assign IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4779 =
	     _theResult_____1__h76814 == 4'd11 && cpReq[37:36] != 2'd2 &&
	     cpReq[9:6] == 4'h9 &&
	     !wci_busy_11 &&
	     wci_respF_11$FULL_N &&
	     !dispatched ;
  assign IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4789 =
	     _theResult_____1__h76814 == 4'd11 && cpReq[37:36] != 2'd2 &&
	     cpReq[9:6] == 4'hA &&
	     !wci_busy_11 &&
	     wci_respF_11$FULL_N &&
	     !dispatched ;
  assign IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4846 =
	     _theResult_____1__h76814 == 4'd12 && cpReq[37:36] != 2'd2 &&
	     cpReq[9:6] == 4'h8 &&
	     !wci_busy_12 &&
	     wci_respF_12$FULL_N &&
	     !dispatched ;
  assign IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4855 =
	     _theResult_____1__h76814 == 4'd12 && cpReq[37:36] != 2'd2 &&
	     cpReq[9:6] == 4'h9 &&
	     !wci_busy_12 &&
	     wci_respF_12$FULL_N &&
	     !dispatched ;
  assign IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4865 =
	     _theResult_____1__h76814 == 4'd12 && cpReq[37:36] != 2'd2 &&
	     cpReq[9:6] == 4'hA &&
	     !wci_busy_12 &&
	     wci_respF_12$FULL_N &&
	     !dispatched ;
  assign IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4922 =
	     _theResult_____1__h76814 == 4'd13 && cpReq[37:36] != 2'd2 &&
	     cpReq[9:6] == 4'h8 &&
	     !wci_busy_13 &&
	     wci_respF_13$FULL_N &&
	     !dispatched ;
  assign IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4931 =
	     _theResult_____1__h76814 == 4'd13 && cpReq[37:36] != 2'd2 &&
	     cpReq[9:6] == 4'h9 &&
	     !wci_busy_13 &&
	     wci_respF_13$FULL_N &&
	     !dispatched ;
  assign IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4941 =
	     _theResult_____1__h76814 == 4'd13 && cpReq[37:36] != 2'd2 &&
	     cpReq[9:6] == 4'hA &&
	     !wci_busy_13 &&
	     wci_respF_13$FULL_N &&
	     !dispatched ;
  assign IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d4998 =
	     _theResult_____1__h76814 == 4'd14 && cpReq[37:36] != 2'd2 &&
	     cpReq[9:6] == 4'h8 &&
	     !wci_busy_14 &&
	     wci_respF_14$FULL_N &&
	     !dispatched ;
  assign IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d5007 =
	     _theResult_____1__h76814 == 4'd14 && cpReq[37:36] != 2'd2 &&
	     cpReq[9:6] == 4'h9 &&
	     !wci_busy_14 &&
	     wci_respF_14$FULL_N &&
	     !dispatched ;
  assign IF_cpReq_363_BITS_37_TO_36_887_EQ_2_888_THEN_c_ETC___d5017 =
	     _theResult_____1__h76814 == 4'd14 && cpReq[37:36] != 2'd2 &&
	     cpReq[9:6] == 4'hA &&
	     !wci_busy_14 &&
	     wci_respF_14$FULL_N &&
	     !dispatched ;
`ifdef not
  assign IF_timeServ_ppsOK_7_THEN_timeServ_ppsExtSync_d_ETC___d5465 =
	     timeServ_ppsOK ?
	       timeServ_ppsExtSync_d2 && !timeServ_ppsExtSyncD :
	       timeServ_delSec != timeServ_fracSeconds[49:48] ;
`endif
  assign IF_wci_lastControlOp_10_713_BIT_3_714_THEN_wci_ETC___d1728 =
	     { wci_lastControlOp_10[3] ? wci_lastControlOp_10[2:0] : 3'b111,
	       wci_lastConfigBE_10[4] ? wci_lastConfigBE_10[3:0] : 4'hF,
	       wci_lastOpWrite_10[1],
	       wci_lastControlOp_10[3],
	       wci_lastConfigBE_10[4],
	       wci_lastConfigAddr_10[32],
	       6'b0,
	       wci_sfCap_10,
	       wci_reqTO_10,
	       wci_reqFAIL_10,
	       wci_reqERR_10 } ;
  assign IF_wci_lastControlOp_11_853_BIT_3_854_THEN_wci_ETC___d1868 =
	     { wci_lastControlOp_11[3] ? wci_lastControlOp_11[2:0] : 3'b111,
	       wci_lastConfigBE_11[4] ? wci_lastConfigBE_11[3:0] : 4'hF,
	       wci_lastOpWrite_11[1],
	       wci_lastControlOp_11[3],
	       wci_lastConfigBE_11[4],
	       wci_lastConfigAddr_11[32],
	       6'b0,
	       wci_sfCap_11,
	       wci_reqTO_11,
	       wci_reqFAIL_11,
	       wci_reqERR_11 } ;
  assign IF_wci_lastControlOp_12_993_BIT_3_994_THEN_wci_ETC___d2008 =
	     { wci_lastControlOp_12[3] ? wci_lastControlOp_12[2:0] : 3'b111,
	       wci_lastConfigBE_12[4] ? wci_lastConfigBE_12[3:0] : 4'hF,
	       wci_lastOpWrite_12[1],
	       wci_lastControlOp_12[3],
	       wci_lastConfigBE_12[4],
	       wci_lastConfigAddr_12[32],
	       6'b0,
	       wci_sfCap_12,
	       wci_reqTO_12,
	       wci_reqFAIL_12,
	       wci_reqERR_12 } ;
  assign IF_wci_lastControlOp_13_133_BIT_3_134_THEN_wci_ETC___d2148 =
	     { wci_lastControlOp_13[3] ? wci_lastControlOp_13[2:0] : 3'b111,
	       wci_lastConfigBE_13[4] ? wci_lastConfigBE_13[3:0] : 4'hF,
	       wci_lastOpWrite_13[1],
	       wci_lastControlOp_13[3],
	       wci_lastConfigBE_13[4],
	       wci_lastConfigAddr_13[32],
	       6'b0,
	       wci_sfCap_13,
	       wci_reqTO_13,
	       wci_reqFAIL_13,
	       wci_reqERR_13 } ;
  assign IF_wci_lastControlOp_13_BIT_3_14_THEN_wci_last_ETC___d328 =
	     { wci_lastControlOp[3] ? wci_lastControlOp[2:0] : 3'b111,
	       wci_lastConfigBE[4] ? wci_lastConfigBE[3:0] : 4'hF,
	       wci_lastOpWrite[1],
	       wci_lastControlOp[3],
	       wci_lastConfigBE[4],
	       wci_lastConfigAddr[32],
	       6'b0,
	       wci_sfCap,
	       wci_reqTO,
	       wci_reqFAIL,
	       wci_reqERR } ;
  assign IF_wci_lastControlOp_14_273_BIT_3_274_THEN_wci_ETC___d2288 =
	     { wci_lastControlOp_14[3] ? wci_lastControlOp_14[2:0] : 3'b111,
	       wci_lastConfigBE_14[4] ? wci_lastConfigBE_14[3:0] : 4'hF,
	       wci_lastOpWrite_14[1],
	       wci_lastControlOp_14[3],
	       wci_lastConfigBE_14[4],
	       wci_lastConfigAddr_14[32],
	       6'b0,
	       wci_sfCap_14,
	       wci_reqTO_14,
	       wci_reqFAIL_14,
	       wci_reqERR_14 } ;
  assign IF_wci_lastControlOp_1_53_BIT_3_54_THEN_wci_la_ETC___d468 =
	     { wci_lastControlOp_1[3] ? wci_lastControlOp_1[2:0] : 3'b111,
	       wci_lastConfigBE_1[4] ? wci_lastConfigBE_1[3:0] : 4'hF,
	       wci_lastOpWrite_1[1],
	       wci_lastControlOp_1[3],
	       wci_lastConfigBE_1[4],
	       wci_lastConfigAddr_1[32],
	       6'b0,
	       wci_sfCap_1,
	       wci_reqTO_1,
	       wci_reqFAIL_1,
	       wci_reqERR_1 } ;
  assign IF_wci_lastControlOp_2_93_BIT_3_94_THEN_wci_la_ETC___d608 =
	     { wci_lastControlOp_2[3] ? wci_lastControlOp_2[2:0] : 3'b111,
	       wci_lastConfigBE_2[4] ? wci_lastConfigBE_2[3:0] : 4'hF,
	       wci_lastOpWrite_2[1],
	       wci_lastControlOp_2[3],
	       wci_lastConfigBE_2[4],
	       wci_lastConfigAddr_2[32],
	       6'b0,
	       wci_sfCap_2,
	       wci_reqTO_2,
	       wci_reqFAIL_2,
	       wci_reqERR_2 } ;
  assign IF_wci_lastControlOp_3_33_BIT_3_34_THEN_wci_la_ETC___d748 =
	     { wci_lastControlOp_3[3] ? wci_lastControlOp_3[2:0] : 3'b111,
	       wci_lastConfigBE_3[4] ? wci_lastConfigBE_3[3:0] : 4'hF,
	       wci_lastOpWrite_3[1],
	       wci_lastControlOp_3[3],
	       wci_lastConfigBE_3[4],
	       wci_lastConfigAddr_3[32],
	       6'b0,
	       wci_sfCap_3,
	       wci_reqTO_3,
	       wci_reqFAIL_3,
	       wci_reqERR_3 } ;
  assign IF_wci_lastControlOp_4_73_BIT_3_74_THEN_wci_la_ETC___d888 =
	     { wci_lastControlOp_4[3] ? wci_lastControlOp_4[2:0] : 3'b111,
	       wci_lastConfigBE_4[4] ? wci_lastConfigBE_4[3:0] : 4'hF,
	       wci_lastOpWrite_4[1],
	       wci_lastControlOp_4[3],
	       wci_lastConfigBE_4[4],
	       wci_lastConfigAddr_4[32],
	       6'b0,
	       wci_sfCap_4,
	       wci_reqTO_4,
	       wci_reqFAIL_4,
	       wci_reqERR_4 } ;
  assign IF_wci_lastControlOp_5_013_BIT_3_014_THEN_wci__ETC___d1028 =
	     { wci_lastControlOp_5[3] ? wci_lastControlOp_5[2:0] : 3'b111,
	       wci_lastConfigBE_5[4] ? wci_lastConfigBE_5[3:0] : 4'hF,
	       wci_lastOpWrite_5[1],
	       wci_lastControlOp_5[3],
	       wci_lastConfigBE_5[4],
	       wci_lastConfigAddr_5[32],
	       6'b0,
	       wci_sfCap_5,
	       wci_reqTO_5,
	       wci_reqFAIL_5,
	       wci_reqERR_5 } ;
  assign IF_wci_lastControlOp_6_153_BIT_3_154_THEN_wci__ETC___d1168 =
	     { wci_lastControlOp_6[3] ? wci_lastControlOp_6[2:0] : 3'b111,
	       wci_lastConfigBE_6[4] ? wci_lastConfigBE_6[3:0] : 4'hF,
	       wci_lastOpWrite_6[1],
	       wci_lastControlOp_6[3],
	       wci_lastConfigBE_6[4],
	       wci_lastConfigAddr_6[32],
	       6'b0,
	       wci_sfCap_6,
	       wci_reqTO_6,
	       wci_reqFAIL_6,
	       wci_reqERR_6 } ;
  assign IF_wci_lastControlOp_7_293_BIT_3_294_THEN_wci__ETC___d1308 =
	     { wci_lastControlOp_7[3] ? wci_lastControlOp_7[2:0] : 3'b111,
	       wci_lastConfigBE_7[4] ? wci_lastConfigBE_7[3:0] : 4'hF,
	       wci_lastOpWrite_7[1],
	       wci_lastControlOp_7[3],
	       wci_lastConfigBE_7[4],
	       wci_lastConfigAddr_7[32],
	       6'b0,
	       wci_sfCap_7,
	       wci_reqTO_7,
	       wci_reqFAIL_7,
	       wci_reqERR_7 } ;
  assign IF_wci_lastControlOp_8_433_BIT_3_434_THEN_wci__ETC___d1448 =
	     { wci_lastControlOp_8[3] ? wci_lastControlOp_8[2:0] : 3'b111,
	       wci_lastConfigBE_8[4] ? wci_lastConfigBE_8[3:0] : 4'hF,
	       wci_lastOpWrite_8[1],
	       wci_lastControlOp_8[3],
	       wci_lastConfigBE_8[4],
	       wci_lastConfigAddr_8[32],
	       6'b0,
	       wci_sfCap_8,
	       wci_reqTO_8,
	       wci_reqFAIL_8,
	       wci_reqERR_8 } ;
  assign IF_wci_lastControlOp_9_573_BIT_3_574_THEN_wci__ETC___d1588 =
	     { wci_lastControlOp_9[3] ? wci_lastControlOp_9[2:0] : 3'b111,
	       wci_lastConfigBE_9[4] ? wci_lastConfigBE_9[3:0] : 4'hF,
	       wci_lastOpWrite_9[1],
	       wci_lastControlOp_9[3],
	       wci_lastConfigBE_9[4],
	       wci_lastConfigAddr_9[32],
	       6'b0,
	       wci_sfCap_9,
	       wci_reqTO_9,
	       wci_reqFAIL_9,
	       wci_reqERR_9 } ;
  assign NOT_cpReq_363_BITS_11_TO_4_366_EQ_0x30_595_649_ETC___d2712 =
	     cpReq[11:4] != 8'h30 && cpReq[11:4] != 8'h34 &&
	     cpReq[11:4] != 8'h38 &&
	     cpReq[11:4] != 8'h3C &&
	     cpReq[11:4] != 8'h40 &&
	     cpReq[11:4] != 8'h44 &&
	     cpReq[11:4] != 8'h48 &&
	     cpReq[11:4] != 8'h4C &&
	     adminResp2F$FULL_N &&
	     !dispatched ;
  assign NOT_cpReq_363_BITS_64_TO_62_364_EQ_0_881_886_A_ETC___d5073 =
	     cpReq[64:62] != 3'd0 && _theResult_____1__h76814 != 4'd0 &&
	     _theResult_____1__h76814 != 4'd1 &&
	     _theResult_____1__h76814 != 4'd2 &&
	     _theResult_____1__h76814 != 4'd3 &&
	     _theResult_____1__h76814 != 4'd4 &&
	     _theResult_____1__h76814 != 4'd5 &&
	     _theResult_____1__h76814 != 4'd6 &&
	     _theResult_____1__h76814 != 4'd7 &&
	     _theResult_____1__h76814 != 4'd8 &&
	     _theResult_____1__h76814 != 4'd9 &&
	     _theResult_____1__h76814 != 4'd10 &&
	     _theResult_____1__h76814 != 4'd11 &&
	     _theResult_____1__h76814 != 4'd12 &&
	     _theResult_____1__h76814 != 4'd13 &&
	     _theResult_____1__h76814 != 4'd14 &&
	     !dispatched ;
  assign NOT_cpReq_363_BITS_64_TO_62_364_EQ_3_877_885_A_ETC___d3976 =
	     cpReq[64:62] != 3'd3 && cpReq[64:62] != 3'd0 &&
	     _theResult_____1__h76814 == 4'd0 &&
	     cpReq[37:36] != 2'd2 &&
	     (cpReq[37:36] != 2'd1 || cpReq[19:9] != 11'd0) &&
	     cpReq[9:6] != 4'h8 &&
	     cpReq[9:6] != 4'h9 &&
	     cpReq[9:6] != 4'hA &&
	     NOT_cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_961_A_ETC___d2962 ;
  assign NOT_cpReq_363_BITS_64_TO_62_364_EQ_3_877_885_A_ETC___d4052 =
	     cpReq[64:62] != 3'd3 && cpReq[64:62] != 3'd0 &&
	     _theResult_____1__h76814 == 4'd1 &&
	     cpReq[37:36] != 2'd2 &&
	     (cpReq[37:36] != 2'd1 || cpReq[19:9] != 11'd0) &&
	     cpReq[9:6] != 4'h8 &&
	     cpReq[9:6] != 4'h9 &&
	     cpReq[9:6] != 4'hA &&
	     NOT_cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_961_A_ETC___d3025 ;
  assign NOT_cpReq_363_BITS_64_TO_62_364_EQ_3_877_885_A_ETC___d4128 =
	     cpReq[64:62] != 3'd3 && cpReq[64:62] != 3'd0 &&
	     _theResult_____1__h76814 == 4'd2 &&
	     cpReq[37:36] != 2'd2 &&
	     (cpReq[37:36] != 2'd1 || cpReq[19:9] != 11'd0) &&
	     cpReq[9:6] != 4'h8 &&
	     cpReq[9:6] != 4'h9 &&
	     cpReq[9:6] != 4'hA &&
	     NOT_cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_961_A_ETC___d3088 ;
  assign NOT_cpReq_363_BITS_64_TO_62_364_EQ_3_877_885_A_ETC___d4204 =
	     cpReq[64:62] != 3'd3 && cpReq[64:62] != 3'd0 &&
	     _theResult_____1__h76814 == 4'd3 &&
	     cpReq[37:36] != 2'd2 &&
	     (cpReq[37:36] != 2'd1 || cpReq[19:9] != 11'd0) &&
	     cpReq[9:6] != 4'h8 &&
	     cpReq[9:6] != 4'h9 &&
	     cpReq[9:6] != 4'hA &&
	     NOT_cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_961_A_ETC___d3151 ;
  assign NOT_cpReq_363_BITS_64_TO_62_364_EQ_3_877_885_A_ETC___d4280 =
	     cpReq[64:62] != 3'd3 && cpReq[64:62] != 3'd0 &&
	     _theResult_____1__h76814 == 4'd4 &&
	     cpReq[37:36] != 2'd2 &&
	     (cpReq[37:36] != 2'd1 || cpReq[19:9] != 11'd0) &&
	     cpReq[9:6] != 4'h8 &&
	     cpReq[9:6] != 4'h9 &&
	     cpReq[9:6] != 4'hA &&
	     NOT_cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_961_A_ETC___d3214 ;
  assign NOT_cpReq_363_BITS_64_TO_62_364_EQ_3_877_885_A_ETC___d4356 =
	     cpReq[64:62] != 3'd3 && cpReq[64:62] != 3'd0 &&
	     _theResult_____1__h76814 == 4'd5 &&
	     cpReq[37:36] != 2'd2 &&
	     (cpReq[37:36] != 2'd1 || cpReq[19:9] != 11'd0) &&
	     cpReq[9:6] != 4'h8 &&
	     cpReq[9:6] != 4'h9 &&
	     cpReq[9:6] != 4'hA &&
	     NOT_cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_961_A_ETC___d3277 ;
  assign NOT_cpReq_363_BITS_64_TO_62_364_EQ_3_877_885_A_ETC___d4432 =
	     cpReq[64:62] != 3'd3 && cpReq[64:62] != 3'd0 &&
	     _theResult_____1__h76814 == 4'd6 &&
	     cpReq[37:36] != 2'd2 &&
	     (cpReq[37:36] != 2'd1 || cpReq[19:9] != 11'd0) &&
	     cpReq[9:6] != 4'h8 &&
	     cpReq[9:6] != 4'h9 &&
	     cpReq[9:6] != 4'hA &&
	     NOT_cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_961_A_ETC___d3340 ;
  assign NOT_cpReq_363_BITS_64_TO_62_364_EQ_3_877_885_A_ETC___d4508 =
	     cpReq[64:62] != 3'd3 && cpReq[64:62] != 3'd0 &&
	     _theResult_____1__h76814 == 4'd7 &&
	     cpReq[37:36] != 2'd2 &&
	     (cpReq[37:36] != 2'd1 || cpReq[19:9] != 11'd0) &&
	     cpReq[9:6] != 4'h8 &&
	     cpReq[9:6] != 4'h9 &&
	     cpReq[9:6] != 4'hA &&
	     NOT_cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_961_A_ETC___d3403 ;
  assign NOT_cpReq_363_BITS_64_TO_62_364_EQ_3_877_885_A_ETC___d4584 =
	     cpReq[64:62] != 3'd3 && cpReq[64:62] != 3'd0 &&
	     _theResult_____1__h76814 == 4'd8 &&
	     cpReq[37:36] != 2'd2 &&
	     (cpReq[37:36] != 2'd1 || cpReq[19:9] != 11'd0) &&
	     cpReq[9:6] != 4'h8 &&
	     cpReq[9:6] != 4'h9 &&
	     cpReq[9:6] != 4'hA &&
	     NOT_cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_961_A_ETC___d3466 ;
  assign NOT_cpReq_363_BITS_64_TO_62_364_EQ_3_877_885_A_ETC___d4660 =
	     cpReq[64:62] != 3'd3 && cpReq[64:62] != 3'd0 &&
	     _theResult_____1__h76814 == 4'd9 &&
	     cpReq[37:36] != 2'd2 &&
	     (cpReq[37:36] != 2'd1 || cpReq[19:9] != 11'd0) &&
	     cpReq[9:6] != 4'h8 &&
	     cpReq[9:6] != 4'h9 &&
	     cpReq[9:6] != 4'hA &&
	     NOT_cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_961_A_ETC___d3529 ;
  assign NOT_cpReq_363_BITS_64_TO_62_364_EQ_3_877_885_A_ETC___d4736 =
	     cpReq[64:62] != 3'd3 && cpReq[64:62] != 3'd0 &&
	     _theResult_____1__h76814 == 4'd10 &&
	     cpReq[37:36] != 2'd2 &&
	     (cpReq[37:36] != 2'd1 || cpReq[19:9] != 11'd0) &&
	     cpReq[9:6] != 4'h8 &&
	     cpReq[9:6] != 4'h9 &&
	     cpReq[9:6] != 4'hA &&
	     NOT_cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_961_A_ETC___d3592 ;
  assign NOT_cpReq_363_BITS_64_TO_62_364_EQ_3_877_885_A_ETC___d4812 =
	     cpReq[64:62] != 3'd3 && cpReq[64:62] != 3'd0 &&
	     _theResult_____1__h76814 == 4'd11 &&
	     cpReq[37:36] != 2'd2 &&
	     (cpReq[37:36] != 2'd1 || cpReq[19:9] != 11'd0) &&
	     cpReq[9:6] != 4'h8 &&
	     cpReq[9:6] != 4'h9 &&
	     cpReq[9:6] != 4'hA &&
	     NOT_cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_961_A_ETC___d3655 ;
  assign NOT_cpReq_363_BITS_64_TO_62_364_EQ_3_877_885_A_ETC___d4888 =
	     cpReq[64:62] != 3'd3 && cpReq[64:62] != 3'd0 &&
	     _theResult_____1__h76814 == 4'd12 &&
	     cpReq[37:36] != 2'd2 &&
	     (cpReq[37:36] != 2'd1 || cpReq[19:9] != 11'd0) &&
	     cpReq[9:6] != 4'h8 &&
	     cpReq[9:6] != 4'h9 &&
	     cpReq[9:6] != 4'hA &&
	     NOT_cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_961_A_ETC___d3718 ;
  assign NOT_cpReq_363_BITS_64_TO_62_364_EQ_3_877_885_A_ETC___d4964 =
	     cpReq[64:62] != 3'd3 && cpReq[64:62] != 3'd0 &&
	     _theResult_____1__h76814 == 4'd13 &&
	     cpReq[37:36] != 2'd2 &&
	     (cpReq[37:36] != 2'd1 || cpReq[19:9] != 11'd0) &&
	     cpReq[9:6] != 4'h8 &&
	     cpReq[9:6] != 4'h9 &&
	     cpReq[9:6] != 4'hA &&
	     NOT_cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_961_A_ETC___d3781 ;
  assign NOT_cpReq_363_BITS_64_TO_62_364_EQ_3_877_885_A_ETC___d5040 =
	     cpReq[64:62] != 3'd3 && cpReq[64:62] != 3'd0 &&
	     _theResult_____1__h76814 == 4'd14 &&
	     cpReq[37:36] != 2'd2 &&
	     (cpReq[37:36] != 2'd1 || cpReq[19:9] != 11'd0) &&
	     cpReq[9:6] != 4'h8 &&
	     cpReq[9:6] != 4'h9 &&
	     cpReq[9:6] != 4'hA &&
	     NOT_cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_961_A_ETC___d3844 ;
  assign NOT_cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_961_A_ETC___d2962 =
	     cpReq[9:6] != 4'hC && !wci_busy && wci_respF$FULL_N &&
	     !dispatched ;
  assign NOT_cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_961_A_ETC___d3025 =
	     cpReq[9:6] != 4'hC && !wci_busy_1 && wci_respF_1$FULL_N &&
	     !dispatched ;
  assign NOT_cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_961_A_ETC___d3088 =
	     cpReq[9:6] != 4'hC && !wci_busy_2 && wci_respF_2$FULL_N &&
	     !dispatched ;
  assign NOT_cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_961_A_ETC___d3151 =
	     cpReq[9:6] != 4'hC && !wci_busy_3 && wci_respF_3$FULL_N &&
	     !dispatched ;
  assign NOT_cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_961_A_ETC___d3214 =
	     cpReq[9:6] != 4'hC && !wci_busy_4 && wci_respF_4$FULL_N &&
	     !dispatched ;
  assign NOT_cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_961_A_ETC___d3277 =
	     cpReq[9:6] != 4'hC && !wci_busy_5 && wci_respF_5$FULL_N &&
	     !dispatched ;
  assign NOT_cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_961_A_ETC___d3340 =
	     cpReq[9:6] != 4'hC && !wci_busy_6 && wci_respF_6$FULL_N &&
	     !dispatched ;
  assign NOT_cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_961_A_ETC___d3403 =
	     cpReq[9:6] != 4'hC && !wci_busy_7 && wci_respF_7$FULL_N &&
	     !dispatched ;
  assign NOT_cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_961_A_ETC___d3466 =
	     cpReq[9:6] != 4'hC && !wci_busy_8 && wci_respF_8$FULL_N &&
	     !dispatched ;
  assign NOT_cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_961_A_ETC___d3529 =
	     cpReq[9:6] != 4'hC && !wci_busy_9 && wci_respF_9$FULL_N &&
	     !dispatched ;
  assign NOT_cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_961_A_ETC___d3592 =
	     cpReq[9:6] != 4'hC && !wci_busy_10 && wci_respF_10$FULL_N &&
	     !dispatched ;
  assign NOT_cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_961_A_ETC___d3655 =
	     cpReq[9:6] != 4'hC && !wci_busy_11 && wci_respF_11$FULL_N &&
	     !dispatched ;
  assign NOT_cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_961_A_ETC___d3718 =
	     cpReq[9:6] != 4'hC && !wci_busy_12 && wci_respF_12$FULL_N &&
	     !dispatched ;
  assign NOT_cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_961_A_ETC___d3781 =
	     cpReq[9:6] != 4'hC && !wci_busy_13 && wci_respF_13$FULL_N &&
	     !dispatched ;
  assign NOT_cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_961_A_ETC___d3844 =
	     cpReq[9:6] != 4'hC && !wci_busy_14 && wci_respF_14$FULL_N &&
	     !dispatched ;
  assign NOT_cpReq_363_BIT_36_924_932_AND_NOT_wci_busy__ETC___d2933 =
	     !cpReq[36] && !wci_busy && wci_respF$FULL_N && !dispatched ;
  assign NOT_cpReq_363_BIT_36_924_932_AND_NOT_wci_busy__ETC___d3000 =
	     !cpReq[36] && !wci_busy_1 && wci_respF_1$FULL_N && !dispatched ;
  assign NOT_cpReq_363_BIT_36_924_932_AND_NOT_wci_busy__ETC___d3063 =
	     !cpReq[36] && !wci_busy_2 && wci_respF_2$FULL_N && !dispatched ;
  assign NOT_cpReq_363_BIT_36_924_932_AND_NOT_wci_busy__ETC___d3126 =
	     !cpReq[36] && !wci_busy_3 && wci_respF_3$FULL_N && !dispatched ;
  assign NOT_cpReq_363_BIT_36_924_932_AND_NOT_wci_busy__ETC___d3189 =
	     !cpReq[36] && !wci_busy_4 && wci_respF_4$FULL_N && !dispatched ;
  assign NOT_cpReq_363_BIT_36_924_932_AND_NOT_wci_busy__ETC___d3252 =
	     !cpReq[36] && !wci_busy_5 && wci_respF_5$FULL_N && !dispatched ;
  assign NOT_cpReq_363_BIT_36_924_932_AND_NOT_wci_busy__ETC___d3315 =
	     !cpReq[36] && !wci_busy_6 && wci_respF_6$FULL_N && !dispatched ;
  assign NOT_cpReq_363_BIT_36_924_932_AND_NOT_wci_busy__ETC___d3378 =
	     !cpReq[36] && !wci_busy_7 && wci_respF_7$FULL_N && !dispatched ;
  assign NOT_cpReq_363_BIT_36_924_932_AND_NOT_wci_busy__ETC___d3441 =
	     !cpReq[36] && !wci_busy_8 && wci_respF_8$FULL_N && !dispatched ;
  assign NOT_cpReq_363_BIT_36_924_932_AND_NOT_wci_busy__ETC___d3504 =
	     !cpReq[36] && !wci_busy_9 && wci_respF_9$FULL_N && !dispatched ;
  assign NOT_cpReq_363_BIT_36_924_932_AND_NOT_wci_busy__ETC___d3567 =
	     !cpReq[36] && !wci_busy_10 && wci_respF_10$FULL_N &&
	     !dispatched ;
  assign NOT_cpReq_363_BIT_36_924_932_AND_NOT_wci_busy__ETC___d3630 =
	     !cpReq[36] && !wci_busy_11 && wci_respF_11$FULL_N &&
	     !dispatched ;
  assign NOT_cpReq_363_BIT_36_924_932_AND_NOT_wci_busy__ETC___d3693 =
	     !cpReq[36] && !wci_busy_12 && wci_respF_12$FULL_N &&
	     !dispatched ;
  assign NOT_cpReq_363_BIT_36_924_932_AND_NOT_wci_busy__ETC___d3756 =
	     !cpReq[36] && !wci_busy_13 && wci_respF_13$FULL_N &&
	     !dispatched ;
  assign NOT_cpReq_363_BIT_36_924_932_AND_NOT_wci_busy__ETC___d3819 =
	     !cpReq[36] && !wci_busy_14 && wci_respF_14$FULL_N &&
	     !dispatched ;
  assign NOT_wci_busy_10_636_536_AND_wci_wReset_n_10_61_ETC___d3549 =
	     !wci_busy_10 && (wci_wReset_n_10 || wci_respF_10$FULL_N) &&
	     !dispatched ;
  assign NOT_wci_busy_11_776_599_AND_wci_wReset_n_11_75_ETC___d3612 =
	     !wci_busy_11 && (wci_wReset_n_11 || wci_respF_11$FULL_N) &&
	     !dispatched ;
  assign NOT_wci_busy_12_916_662_AND_wci_wReset_n_12_89_ETC___d3675 =
	     !wci_busy_12 && (wci_wReset_n_12 || wci_respF_12$FULL_N) &&
	     !dispatched ;
  assign NOT_wci_busy_13_056_725_AND_wci_wReset_n_13_03_ETC___d3738 =
	     !wci_busy_13 && (wci_wReset_n_13 || wci_respF_13$FULL_N) &&
	     !dispatched ;
  assign NOT_wci_busy_14_196_788_AND_wci_wReset_n_14_17_ETC___d3801 =
	     !wci_busy_14 && (wci_wReset_n_14 || wci_respF_14$FULL_N) &&
	     !dispatched ;
  assign NOT_wci_busy_1_76_969_AND_wci_wReset_n_1_56_OR_ETC___d2982 =
	     !wci_busy_1 && (wci_wReset_n_1 || wci_respF_1$FULL_N) &&
	     !dispatched ;
  assign NOT_wci_busy_2_16_032_AND_wci_wReset_n_2_96_OR_ETC___d3045 =
	     !wci_busy_2 && (wci_wReset_n_2 || wci_respF_2$FULL_N) &&
	     !dispatched ;
  assign NOT_wci_busy_36_886_AND_wci_wReset_n_16_OR_wci_ETC___d2904 =
	     !wci_busy && (wci_wReset_n || wci_respF$FULL_N) && !dispatched ;
  assign NOT_wci_busy_3_56_095_AND_wci_wReset_n_3_36_OR_ETC___d3108 =
	     !wci_busy_3 && (wci_wReset_n_3 || wci_respF_3$FULL_N) &&
	     !dispatched ;
  assign NOT_wci_busy_4_96_158_AND_wci_wReset_n_4_76_OR_ETC___d3171 =
	     !wci_busy_4 && (wci_wReset_n_4 || wci_respF_4$FULL_N) &&
	     !dispatched ;
  assign NOT_wci_busy_5_36_221_AND_wci_wReset_n_5_16_OR_ETC___d3234 =
	     !wci_busy_5 && (wci_wReset_n_5 || wci_respF_5$FULL_N) &&
	     !dispatched ;
  assign NOT_wci_busy_6_076_284_AND_wci_wReset_n_6_056__ETC___d3297 =
	     !wci_busy_6 && (wci_wReset_n_6 || wci_respF_6$FULL_N) &&
	     !dispatched ;
  assign NOT_wci_busy_7_216_347_AND_wci_wReset_n_7_196__ETC___d3360 =
	     !wci_busy_7 && (wci_wReset_n_7 || wci_respF_7$FULL_N) &&
	     !dispatched ;
  assign NOT_wci_busy_8_356_410_AND_wci_wReset_n_8_336__ETC___d3423 =
	     !wci_busy_8 && (wci_wReset_n_8 || wci_respF_8$FULL_N) &&
	     !dispatched ;
  assign NOT_wci_busy_9_496_473_AND_wci_wReset_n_9_476__ETC___d3486 =
	     !wci_busy_9 && (wci_wReset_n_9 || wci_respF_9$FULL_N) &&
	     !dispatched ;
`ifdef not
  assign _281474976710656_MINUS_timeServ_delSecond_BITS__ETC__q2 =
	     _281474976710656_MINUS_timeServ_delSecond__q1[49:28] ;
  assign _281474976710656_MINUS_timeServ_delSecond__q1 =
	     50'h1000000000000 - timeServ_delSecond ;
`endif
  assign _theResult_____1__h76796 =
	     (cpReq[61:60] == 2'd2) ? wn___1__h77585 : wn__h76795 ;
  assign _theResult_____1__h76814 =
	     (cpReq[37:36] == 2'd2) ? wn___1__h77585 : wn__h76795 ;
  assign bAddr__h113843 = { cpReqF$D_OUT[57:36], 2'b0 } ;
  assign bAddr__h114303 = { cpReqF$D_OUT[25:4], 2'b0 } ;
  assign cpReq_363_BITS_11_TO_4_366_EQ_0x30_595_OR_cpRe_ETC___d2632 =
	     (cpReq[11:4] == 8'h30 || cpReq[11:4] == 8'h34 ||
	      cpReq[11:4] == 8'h38 ||
	      cpReq[11:4] == 8'h3C ||
	      cpReq[11:4] == 8'h40 ||
	      cpReq[11:4] == 8'h44 ||
	      cpReq[11:4] == 8'h48) &&
	     adminResp2F$FULL_N &&
	     !dispatched ;
  assign cpReq_363_BITS_11_TO_4_366_ULT_0x30___d2438 = cpReq[11:4] < 8'h30 ;
  assign cpReq_363_BITS_11_TO_4_366_ULT_0xC0___d2594 = cpReq[11:4] < 8'hC0 ;
  assign cpReq_363_BITS_27_TO_4_436_ULT_0x1000___d2866 =
	     cpReq[27:4] < 24'h001000 ;
  assign cpReq_363_BITS_27_TO_4_436_ULT_0x100___d2437 =
	     cpReq[27:4] < 24'h000100 ;
  assign cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_AND_NOT_w_ETC___d2953 =
	     cpReq[9:6] == 4'hC && !wci_busy && wci_respF$FULL_N &&
	     !dispatched ;
  assign cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_AND_NOT_w_ETC___d3019 =
	     cpReq[9:6] == 4'hC && !wci_busy_1 && wci_respF_1$FULL_N &&
	     !dispatched ;
  assign cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_AND_NOT_w_ETC___d3082 =
	     cpReq[9:6] == 4'hC && !wci_busy_2 && wci_respF_2$FULL_N &&
	     !dispatched ;
  assign cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_AND_NOT_w_ETC___d3145 =
	     cpReq[9:6] == 4'hC && !wci_busy_3 && wci_respF_3$FULL_N &&
	     !dispatched ;
  assign cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_AND_NOT_w_ETC___d3208 =
	     cpReq[9:6] == 4'hC && !wci_busy_4 && wci_respF_4$FULL_N &&
	     !dispatched ;
  assign cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_AND_NOT_w_ETC___d3271 =
	     cpReq[9:6] == 4'hC && !wci_busy_5 && wci_respF_5$FULL_N &&
	     !dispatched ;
  assign cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_AND_NOT_w_ETC___d3334 =
	     cpReq[9:6] == 4'hC && !wci_busy_6 && wci_respF_6$FULL_N &&
	     !dispatched ;
  assign cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_AND_NOT_w_ETC___d3397 =
	     cpReq[9:6] == 4'hC && !wci_busy_7 && wci_respF_7$FULL_N &&
	     !dispatched ;
  assign cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_AND_NOT_w_ETC___d3460 =
	     cpReq[9:6] == 4'hC && !wci_busy_8 && wci_respF_8$FULL_N &&
	     !dispatched ;
  assign cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_AND_NOT_w_ETC___d3523 =
	     cpReq[9:6] == 4'hC && !wci_busy_9 && wci_respF_9$FULL_N &&
	     !dispatched ;
  assign cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_AND_NOT_w_ETC___d3586 =
	     cpReq[9:6] == 4'hC && !wci_busy_10 && wci_respF_10$FULL_N &&
	     !dispatched ;
  assign cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_AND_NOT_w_ETC___d3649 =
	     cpReq[9:6] == 4'hC && !wci_busy_11 && wci_respF_11$FULL_N &&
	     !dispatched ;
  assign cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_AND_NOT_w_ETC___d3712 =
	     cpReq[9:6] == 4'hC && !wci_busy_12 && wci_respF_12$FULL_N &&
	     !dispatched ;
  assign cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_AND_NOT_w_ETC___d3775 =
	     cpReq[9:6] == 4'hC && !wci_busy_13 && wci_respF_13$FULL_N &&
	     !dispatched ;
  assign cpReq_363_BITS_9_TO_6_796_EQ_0xC_835_AND_NOT_w_ETC___d3838 =
	     cpReq[9:6] == 4'hC && !wci_busy_14 && wci_respF_14$FULL_N &&
	     !dispatched ;
  assign cpReq_363_BIT_36_924_AND_NOT_wci_busy_10_636_5_ETC___d3560 =
	     cpReq[36] && !wci_busy_10 && wci_respF_10$FULL_N && !dispatched ;
  assign cpReq_363_BIT_36_924_AND_NOT_wci_busy_11_776_5_ETC___d3623 =
	     cpReq[36] && !wci_busy_11 && wci_respF_11$FULL_N && !dispatched ;
  assign cpReq_363_BIT_36_924_AND_NOT_wci_busy_12_916_6_ETC___d3686 =
	     cpReq[36] && !wci_busy_12 && wci_respF_12$FULL_N && !dispatched ;
  assign cpReq_363_BIT_36_924_AND_NOT_wci_busy_13_056_7_ETC___d3749 =
	     cpReq[36] && !wci_busy_13 && wci_respF_13$FULL_N && !dispatched ;
  assign cpReq_363_BIT_36_924_AND_NOT_wci_busy_14_196_7_ETC___d3812 =
	     cpReq[36] && !wci_busy_14 && wci_respF_14$FULL_N && !dispatched ;
  assign cpReq_363_BIT_36_924_AND_NOT_wci_busy_1_76_969_ETC___d2993 =
	     cpReq[36] && !wci_busy_1 && wci_respF_1$FULL_N && !dispatched ;
  assign cpReq_363_BIT_36_924_AND_NOT_wci_busy_2_16_032_ETC___d3056 =
	     cpReq[36] && !wci_busy_2 && wci_respF_2$FULL_N && !dispatched ;
  assign cpReq_363_BIT_36_924_AND_NOT_wci_busy_36_886_A_ETC___d2925 =
	     cpReq[36] && !wci_busy && wci_respF$FULL_N && !dispatched ;
  assign cpReq_363_BIT_36_924_AND_NOT_wci_busy_3_56_095_ETC___d3119 =
	     cpReq[36] && !wci_busy_3 && wci_respF_3$FULL_N && !dispatched ;
  assign cpReq_363_BIT_36_924_AND_NOT_wci_busy_4_96_158_ETC___d3182 =
	     cpReq[36] && !wci_busy_4 && wci_respF_4$FULL_N && !dispatched ;
  assign cpReq_363_BIT_36_924_AND_NOT_wci_busy_5_36_221_ETC___d3245 =
	     cpReq[36] && !wci_busy_5 && wci_respF_5$FULL_N && !dispatched ;
  assign cpReq_363_BIT_36_924_AND_NOT_wci_busy_6_076_28_ETC___d3308 =
	     cpReq[36] && !wci_busy_6 && wci_respF_6$FULL_N && !dispatched ;
  assign cpReq_363_BIT_36_924_AND_NOT_wci_busy_7_216_34_ETC___d3371 =
	     cpReq[36] && !wci_busy_7 && wci_respF_7$FULL_N && !dispatched ;
  assign cpReq_363_BIT_36_924_AND_NOT_wci_busy_8_356_41_ETC___d3434 =
	     cpReq[36] && !wci_busy_8 && wci_respF_8$FULL_N && !dispatched ;
  assign cpReq_363_BIT_36_924_AND_NOT_wci_busy_9_496_47_ETC___d3497 =
	     cpReq[36] && !wci_busy_9 && wci_respF_9$FULL_N && !dispatched ;
  assign cpStatus__h75932 = { 28'd0, rogueTLP } ;
  assign crr_data__h76602 =
	     adminRespF$D_OUT[32] ? adminRespF$D_OUT[31:0] : 32'hDEADC0DE ;
`ifdef not
  assign rom_serverAdapter_cnt_29_PLUS_IF_rom_serverAda_ETC___d135 =
	     rom_serverAdapter_cnt +
	     (WILL_FIRE_RL_rom_serverAdapter_stageReadResponseAlways ?
		3'd1 :
		3'd0) +
	     (rom_serverAdapter_outData_deqCalled$whas ? 3'd7 : 3'd0) ;
  assign timeServ_ppsExtSync_d2_2_AND_NOT_timeServ_ppsE_ETC___d61 =
	     timeServ_ppsExtSync_d2 && !timeServ_ppsExtSyncD &&
	     (timeServ_refFromRise_3_ULE_199800000___d5459 ||
	      !timeServ_refFromRise_3_ULT_200200000___d5878) ||
	     timeServ_refFromRise > 28'd200200000 ;
  assign timeServ_ppsExtSync_d2_2_AND_NOT_timeServ_ppsE_ETC___d70 =
	     timeServ_ppsExtSync_d2 && !timeServ_ppsExtSyncD &&
	     !timeServ_refFromRise_3_ULE_199800000___d5459 &&
	     timeServ_refFromRise_3_ULT_200200000___d5878 &&
	     timeServ_ppsOK &&
	     !timeServ_disableServo$dD_OUT ;
  assign timeServ_refFromRise_3_ULE_199800000___d5459 =
	     timeServ_refFromRise <= 28'd199800000 ;
  assign timeServ_refFromRise_3_ULT_200200000___d5878 =
	     timeServ_refFromRise < 28'd200200000 ;
`endif
  assign toCount__h11764 = 32'd1 << wci_wTimeout ;
  assign toCount__h16210 = 32'd1 << wci_wTimeout_1 ;
  assign toCount__h20650 = 32'd1 << wci_wTimeout_2 ;
  assign toCount__h25090 = 32'd1 << wci_wTimeout_3 ;
  assign toCount__h29530 = 32'd1 << wci_wTimeout_4 ;
  assign toCount__h33970 = 32'd1 << wci_wTimeout_5 ;
  assign toCount__h38410 = 32'd1 << wci_wTimeout_6 ;
  assign toCount__h42850 = 32'd1 << wci_wTimeout_7 ;
  assign toCount__h47290 = 32'd1 << wci_wTimeout_8 ;
  assign toCount__h51730 = 32'd1 << wci_wTimeout_9 ;
  assign toCount__h56170 = 32'd1 << wci_wTimeout_10 ;
  assign toCount__h60610 = 32'd1 << wci_wTimeout_11 ;
  assign toCount__h65050 = 32'd1 << wci_wTimeout_12 ;
  assign toCount__h69490 = 32'd1 << wci_wTimeout_13 ;
  assign toCount__h73930 = 32'd1 << wci_wTimeout_14 ;
  assign wciAddr__h78327 = { wci_pageWindow, cpReq[23:4] } ;
  assign wciAddr__h78395 = { wci_pageWindow_1, cpReq[23:4] } ;
  assign wciAddr__h78461 = { wci_pageWindow_2, cpReq[23:4] } ;
  assign wciAddr__h78527 = { wci_pageWindow_3, cpReq[23:4] } ;
  assign wciAddr__h78593 = { wci_pageWindow_4, cpReq[23:4] } ;
  assign wciAddr__h78659 = { wci_pageWindow_5, cpReq[23:4] } ;
  assign wciAddr__h78725 = { wci_pageWindow_6, cpReq[23:4] } ;
  assign wciAddr__h78791 = { wci_pageWindow_7, cpReq[23:4] } ;
  assign wciAddr__h78857 = { wci_pageWindow_8, cpReq[23:4] } ;
  assign wciAddr__h78923 = { wci_pageWindow_9, cpReq[23:4] } ;
  assign wciAddr__h78989 = { wci_pageWindow_10, cpReq[23:4] } ;
  assign wciAddr__h79055 = { wci_pageWindow_11, cpReq[23:4] } ;
  assign wciAddr__h79121 = { wci_pageWindow_12, cpReq[23:4] } ;
  assign wciAddr__h79187 = { wci_pageWindow_13, cpReq[23:4] } ;
  assign wciAddr__h79253 = { wci_pageWindow_14, cpReq[23:4] } ;
  assign wci_respTimr_10_628_ULT_1_SL_wci_wTimeout_10_6_ETC___d5889 =
	     wci_respTimr_10 < toCount__h56170 ;
  assign wci_respTimr_11_768_ULT_1_SL_wci_wTimeout_11_7_ETC___d5890 =
	     wci_respTimr_11 < toCount__h60610 ;
  assign wci_respTimr_12_908_ULT_1_SL_wci_wTimeout_12_9_ETC___d5891 =
	     wci_respTimr_12 < toCount__h65050 ;
  assign wci_respTimr_13_048_ULT_1_SL_wci_wTimeout_13_0_ETC___d5892 =
	     wci_respTimr_13 < toCount__h69490 ;
  assign wci_respTimr_14_188_ULT_1_SL_wci_wTimeout_14_1_ETC___d5893 =
	     wci_respTimr_14 < toCount__h73930 ;
  assign wci_respTimr_1_68_ULT_1_SL_wci_wTimeout_1_69_70___d5880 =
	     wci_respTimr_1 < toCount__h16210 ;
  assign wci_respTimr_28_ULT_1_SL_wci_wTimeout_29_30___d5879 =
	     wci_respTimr < toCount__h11764 ;
  assign wci_respTimr_2_08_ULT_1_SL_wci_wTimeout_2_09_10___d5881 =
	     wci_respTimr_2 < toCount__h20650 ;
  assign wci_respTimr_3_48_ULT_1_SL_wci_wTimeout_3_49_50___d5882 =
	     wci_respTimr_3 < toCount__h25090 ;
  assign wci_respTimr_4_88_ULT_1_SL_wci_wTimeout_4_89_90___d5883 =
	     wci_respTimr_4 < toCount__h29530 ;
  assign wci_respTimr_5_28_ULT_1_SL_wci_wTimeout_5_29_30___d5884 =
	     wci_respTimr_5 < toCount__h33970 ;
  assign wci_respTimr_6_068_ULT_1_SL_wci_wTimeout_6_069_ETC___d5885 =
	     wci_respTimr_6 < toCount__h38410 ;
  assign wci_respTimr_7_208_ULT_1_SL_wci_wTimeout_7_209_ETC___d5886 =
	     wci_respTimr_7 < toCount__h42850 ;
  assign wci_respTimr_8_348_ULT_1_SL_wci_wTimeout_8_349_ETC___d5887 =
	     wci_respTimr_8 < toCount__h47290 ;
  assign wci_respTimr_9_488_ULT_1_SL_wci_wTimeout_9_489_ETC___d5888 =
	     wci_respTimr_9 < toCount__h51730 ;
  assign wci_wReset_n_10_616_AND_NOT_wci_busy_10_636_53_ETC___d3539 =
	     wci_wReset_n_10 && !wci_busy_10 && !wci_reqF_10_c_r &&
	     !dispatched ;
  assign wci_wReset_n_11_756_AND_NOT_wci_busy_11_776_59_ETC___d3602 =
	     wci_wReset_n_11 && !wci_busy_11 && !wci_reqF_11_c_r &&
	     !dispatched ;
  assign wci_wReset_n_12_896_AND_NOT_wci_busy_12_916_66_ETC___d3665 =
	     wci_wReset_n_12 && !wci_busy_12 && !wci_reqF_12_c_r &&
	     !dispatched ;
  assign wci_wReset_n_13_036_AND_NOT_wci_busy_13_056_72_ETC___d3728 =
	     wci_wReset_n_13 && !wci_busy_13 && !wci_reqF_13_c_r &&
	     !dispatched ;
  assign wci_wReset_n_14_176_AND_NOT_wci_busy_14_196_78_ETC___d3791 =
	     wci_wReset_n_14 && !wci_busy_14 && !wci_reqF_14_c_r &&
	     !dispatched ;
  assign wci_wReset_n_16_AND_NOT_wci_busy_36_886_AND_NO_ETC___d2889 =
	     wci_wReset_n && !wci_busy && !wci_reqF_c_r && !dispatched ;
  assign wci_wReset_n_1_56_AND_NOT_wci_busy_1_76_969_AN_ETC___d2972 =
	     wci_wReset_n_1 && !wci_busy_1 && !wci_reqF_1_c_r && !dispatched ;
  assign wci_wReset_n_2_96_AND_NOT_wci_busy_2_16_032_AN_ETC___d3035 =
	     wci_wReset_n_2 && !wci_busy_2 && !wci_reqF_2_c_r && !dispatched ;
  assign wci_wReset_n_3_36_AND_NOT_wci_busy_3_56_095_AN_ETC___d3098 =
	     wci_wReset_n_3 && !wci_busy_3 && !wci_reqF_3_c_r && !dispatched ;
  assign wci_wReset_n_4_76_AND_NOT_wci_busy_4_96_158_AN_ETC___d3161 =
	     wci_wReset_n_4 && !wci_busy_4 && !wci_reqF_4_c_r && !dispatched ;
  assign wci_wReset_n_5_16_AND_NOT_wci_busy_5_36_221_AN_ETC___d3224 =
	     wci_wReset_n_5 && !wci_busy_5 && !wci_reqF_5_c_r && !dispatched ;
  assign wci_wReset_n_6_056_AND_NOT_wci_busy_6_076_284__ETC___d3287 =
	     wci_wReset_n_6 && !wci_busy_6 && !wci_reqF_6_c_r && !dispatched ;
  assign wci_wReset_n_7_196_AND_NOT_wci_busy_7_216_347__ETC___d3350 =
	     wci_wReset_n_7 && !wci_busy_7 && !wci_reqF_7_c_r && !dispatched ;
  assign wci_wReset_n_8_336_AND_NOT_wci_busy_8_356_410__ETC___d3413 =
	     wci_wReset_n_8 && !wci_busy_8 && !wci_reqF_8_c_r && !dispatched ;
  assign wci_wReset_n_9_476_AND_NOT_wci_busy_9_496_473__ETC___d3476 =
	     wci_wReset_n_9 && !wci_busy_9 && !wci_reqF_9_c_r && !dispatched ;
  assign wci_wciResponse_10_wget__623_BITS_33_TO_32_624_ETC___d1652 =
	     wci_wciResponse_10$wget[33:32] == 2'd0 &&
	     !wci_respTimr_10_628_ULT_1_SL_wci_wTimeout_10_6_ETC___d5889 &&
	     (wci_reqPend_10 == 2'd1 || wci_reqPend_10 == 2'd2 ||
	      wci_reqPend_10 == 2'd3) ;
  assign wci_wciResponse_11_wget__763_BITS_33_TO_32_764_ETC___d1792 =
	     wci_wciResponse_11$wget[33:32] == 2'd0 &&
	     !wci_respTimr_11_768_ULT_1_SL_wci_wTimeout_11_7_ETC___d5890 &&
	     (wci_reqPend_11 == 2'd1 || wci_reqPend_11 == 2'd2 ||
	      wci_reqPend_11 == 2'd3) ;
  assign wci_wciResponse_12_wget__903_BITS_33_TO_32_904_ETC___d1932 =
	     wci_wciResponse_12$wget[33:32] == 2'd0 &&
	     !wci_respTimr_12_908_ULT_1_SL_wci_wTimeout_12_9_ETC___d5891 &&
	     (wci_reqPend_12 == 2'd1 || wci_reqPend_12 == 2'd2 ||
	      wci_reqPend_12 == 2'd3) ;
  assign wci_wciResponse_13_wget__043_BITS_33_TO_32_044_ETC___d2072 =
	     wci_wciResponse_13$wget[33:32] == 2'd0 &&
	     !wci_respTimr_13_048_ULT_1_SL_wci_wTimeout_13_0_ETC___d5892 &&
	     (wci_reqPend_13 == 2'd1 || wci_reqPend_13 == 2'd2 ||
	      wci_reqPend_13 == 2'd3) ;
  assign wci_wciResponse_14_wget__183_BITS_33_TO_32_184_ETC___d2212 =
	     wci_wciResponse_14$wget[33:32] == 2'd0 &&
	     !wci_respTimr_14_188_ULT_1_SL_wci_wTimeout_14_1_ETC___d5893 &&
	     (wci_reqPend_14 == 2'd1 || wci_reqPend_14 == 2'd2 ||
	      wci_reqPend_14 == 2'd3) ;
  assign wci_wciResponse_1_wget__63_BITS_33_TO_32_64_EQ_ETC___d392 =
	     wci_wciResponse_1$wget[33:32] == 2'd0 &&
	     !wci_respTimr_1_68_ULT_1_SL_wci_wTimeout_1_69_70___d5880 &&
	     (wci_reqPend_1 == 2'd1 || wci_reqPend_1 == 2'd2 ||
	      wci_reqPend_1 == 2'd3) ;
  assign wci_wciResponse_2_wget__03_BITS_33_TO_32_04_EQ_ETC___d532 =
	     wci_wciResponse_2$wget[33:32] == 2'd0 &&
	     !wci_respTimr_2_08_ULT_1_SL_wci_wTimeout_2_09_10___d5881 &&
	     (wci_reqPend_2 == 2'd1 || wci_reqPend_2 == 2'd2 ||
	      wci_reqPend_2 == 2'd3) ;
  assign wci_wciResponse_3_wget__43_BITS_33_TO_32_44_EQ_ETC___d672 =
	     wci_wciResponse_3$wget[33:32] == 2'd0 &&
	     !wci_respTimr_3_48_ULT_1_SL_wci_wTimeout_3_49_50___d5882 &&
	     (wci_reqPend_3 == 2'd1 || wci_reqPend_3 == 2'd2 ||
	      wci_reqPend_3 == 2'd3) ;
  assign wci_wciResponse_4_wget__83_BITS_33_TO_32_84_EQ_ETC___d812 =
	     wci_wciResponse_4$wget[33:32] == 2'd0 &&
	     !wci_respTimr_4_88_ULT_1_SL_wci_wTimeout_4_89_90___d5883 &&
	     (wci_reqPend_4 == 2'd1 || wci_reqPend_4 == 2'd2 ||
	      wci_reqPend_4 == 2'd3) ;
  assign wci_wciResponse_5_wget__23_BITS_33_TO_32_24_EQ_ETC___d952 =
	     wci_wciResponse_5$wget[33:32] == 2'd0 &&
	     !wci_respTimr_5_28_ULT_1_SL_wci_wTimeout_5_29_30___d5884 &&
	     (wci_reqPend_5 == 2'd1 || wci_reqPend_5 == 2'd2 ||
	      wci_reqPend_5 == 2'd3) ;
  assign wci_wciResponse_6_wget__063_BITS_33_TO_32_064__ETC___d1092 =
	     wci_wciResponse_6$wget[33:32] == 2'd0 &&
	     !wci_respTimr_6_068_ULT_1_SL_wci_wTimeout_6_069_ETC___d5885 &&
	     (wci_reqPend_6 == 2'd1 || wci_reqPend_6 == 2'd2 ||
	      wci_reqPend_6 == 2'd3) ;
  assign wci_wciResponse_7_wget__203_BITS_33_TO_32_204__ETC___d1232 =
	     wci_wciResponse_7$wget[33:32] == 2'd0 &&
	     !wci_respTimr_7_208_ULT_1_SL_wci_wTimeout_7_209_ETC___d5886 &&
	     (wci_reqPend_7 == 2'd1 || wci_reqPend_7 == 2'd2 ||
	      wci_reqPend_7 == 2'd3) ;
  assign wci_wciResponse_8_wget__343_BITS_33_TO_32_344__ETC___d1372 =
	     wci_wciResponse_8$wget[33:32] == 2'd0 &&
	     !wci_respTimr_8_348_ULT_1_SL_wci_wTimeout_8_349_ETC___d5887 &&
	     (wci_reqPend_8 == 2'd1 || wci_reqPend_8 == 2'd2 ||
	      wci_reqPend_8 == 2'd3) ;
  assign wci_wciResponse_9_wget__483_BITS_33_TO_32_484__ETC___d1512 =
	     wci_wciResponse_9$wget[33:32] == 2'd0 &&
	     !wci_respTimr_9_488_ULT_1_SL_wci_wTimeout_9_489_ETC___d5888 &&
	     (wci_reqPend_9 == 2'd1 || wci_reqPend_9 == 2'd2 ||
	      wci_reqPend_9 == 2'd3) ;
  assign wci_wciResponse_wget__23_BITS_33_TO_32_24_EQ_0_ETC___d252 =
	     wci_wciResponse$wget[33:32] == 2'd0 &&
	     !wci_respTimr_28_ULT_1_SL_wci_wTimeout_29_30___d5879 &&
	     (wci_reqPend == 2'd1 || wci_reqPend == 2'd2 ||
	      wci_reqPend == 2'd3) ;
  assign wn___1__h77585 = cpReq[27:24] - 4'd1 ;
  assign wn__h76795 = cpReq[23:20] - 4'd1 ;
  assign x__h106341 =
	     { wci_slvPresent_14,
	       wci_slvPresent_13,
	       wci_slvPresent_12,
	       wci_slvPresent_11,
	       wci_slvPresent_10,
	       wci_slvPresent_9,
	       wci_slvPresent_8,
	       wci_slvPresent_7,
	       wci_slvPresent_6,
	       wci_slvPresent_5,
	       wci_slvPresent_4,
	       wci_slvPresent_3,
	       wci_slvPresent_2,
	       wci_slvPresent_1,
	       wci_slvPresent } ;
  assign x__h106890 =
	     { wci_wStatus_14[15:0] != 16'd0,
	       wci_wStatus_13[15:0] != 16'd0,
	       wci_wStatus_12[15:0] != 16'd0,
	       wci_wStatus_11[15:0] != 16'd0,
	       wci_wStatus_10[15:0] != 16'd0,
	       wci_wStatus_9[15:0] != 16'd0,
	       wci_wStatus_8[15:0] != 16'd0,
	       wci_wStatus_7[15:0] != 16'd0,
	       wci_wStatus_6[15:0] != 16'd0,
	       wci_wStatus_5[15:0] != 16'd0,
	       wci_wStatus_4[15:0] != 16'd0,
	       wci_wStatus_3[15:0] != 16'd0,
	       wci_wStatus_2[15:0] != 16'd0,
	       wci_wStatus_1[15:0] != 16'd0,
	       wci_wStatus[15:0] != 16'd0 } ;
  assign x__h11924 = wci_respTimr + 32'd1 ;
  assign x__h16367 = wci_respTimr_1 + 32'd1 ;
  assign x__h20807 = wci_respTimr_2 + 32'd1 ;
  assign x__h25247 = wci_respTimr_3 + 32'd1 ;
  assign x__h29687 = wci_respTimr_4 + 32'd1 ;
  assign x__h34127 = wci_respTimr_5 + 32'd1 ;
`ifdef not
  assign x__h3700 = { 2'b0, x_f__h4848 } ;
`endif
  assign x__h38567 = wci_respTimr_6 + 32'd1 ;
  assign x__h43007 = wci_respTimr_7 + 32'd1 ;
`ifdef not
  assign x__h4421 =
	     { {28{_281474976710656_MINUS_timeServ_delSecond_BITS__ETC__q2[21]}},
	       _281474976710656_MINUS_timeServ_delSecond_BITS__ETC__q2 } ;
  assign x__h4649 = timeServ_fracSeconds + timeServ_fracInc ;
  assign x__h4715 = timeServ_refSecCount + 32'd1 ;
`endif
  assign x__h47447 = wci_respTimr_8 + 32'd1 ;
  assign x__h51887 = wci_respTimr_9 + 32'd1 ;
  assign x__h56327 = wci_respTimr_10 + 32'd1 ;
  assign x__h60767 = wci_respTimr_11 + 32'd1 ;
  assign x__h65207 = wci_respTimr_12 + 32'd1 ;
  assign x__h69647 = wci_respTimr_13 + 32'd1 ;
  assign x__h74087 = wci_respTimr_14 + 32'd1 ;
  assign x__h98553 = { cpReq[8:6], 2'b0 } ;
  assign x_addr__h98551 = { 27'd0, x__h98553 } ;
  assign x_data__h104757 = { wci_wReset_n, 26'd0, wci_wTimeout } ;
  assign x_data__h104763 =
	     wci_lastConfigAddr[32] ?
	       wci_lastConfigAddr[31:0] :
	       32'hFFFFFFFF ;
  assign x_data__h104810 = { wci_wReset_n_1, 26'd0, wci_wTimeout_1 } ;
  assign x_data__h104816 =
	     wci_lastConfigAddr_1[32] ?
	       wci_lastConfigAddr_1[31:0] :
	       32'hFFFFFFFF ;
  assign x_data__h104863 = { wci_wReset_n_2, 26'd0, wci_wTimeout_2 } ;
  assign x_data__h104869 =
	     wci_lastConfigAddr_2[32] ?
	       wci_lastConfigAddr_2[31:0] :
	       32'hFFFFFFFF ;
  assign x_data__h104916 = { wci_wReset_n_3, 26'd0, wci_wTimeout_3 } ;
  assign x_data__h104922 =
	     wci_lastConfigAddr_3[32] ?
	       wci_lastConfigAddr_3[31:0] :
	       32'hFFFFFFFF ;
  assign x_data__h104969 = { wci_wReset_n_4, 26'd0, wci_wTimeout_4 } ;
  assign x_data__h104975 =
	     wci_lastConfigAddr_4[32] ?
	       wci_lastConfigAddr_4[31:0] :
	       32'hFFFFFFFF ;
  assign x_data__h105022 = { wci_wReset_n_5, 26'd0, wci_wTimeout_5 } ;
  assign x_data__h105028 =
	     wci_lastConfigAddr_5[32] ?
	       wci_lastConfigAddr_5[31:0] :
	       32'hFFFFFFFF ;
  assign x_data__h105075 = { wci_wReset_n_6, 26'd0, wci_wTimeout_6 } ;
  assign x_data__h105081 =
	     wci_lastConfigAddr_6[32] ?
	       wci_lastConfigAddr_6[31:0] :
	       32'hFFFFFFFF ;
  assign x_data__h105128 = { wci_wReset_n_7, 26'd0, wci_wTimeout_7 } ;
  assign x_data__h105134 =
	     wci_lastConfigAddr_7[32] ?
	       wci_lastConfigAddr_7[31:0] :
	       32'hFFFFFFFF ;
  assign x_data__h105181 = { wci_wReset_n_8, 26'd0, wci_wTimeout_8 } ;
  assign x_data__h105187 =
	     wci_lastConfigAddr_8[32] ?
	       wci_lastConfigAddr_8[31:0] :
	       32'hFFFFFFFF ;
  assign x_data__h105234 = { wci_wReset_n_9, 26'd0, wci_wTimeout_9 } ;
  assign x_data__h105240 =
	     wci_lastConfigAddr_9[32] ?
	       wci_lastConfigAddr_9[31:0] :
	       32'hFFFFFFFF ;
  assign x_data__h105287 = { wci_wReset_n_10, 26'd0, wci_wTimeout_10 } ;
  assign x_data__h105293 =
	     wci_lastConfigAddr_10[32] ?
	       wci_lastConfigAddr_10[31:0] :
	       32'hFFFFFFFF ;
  assign x_data__h105340 = { wci_wReset_n_11, 26'd0, wci_wTimeout_11 } ;
  assign x_data__h105346 =
	     wci_lastConfigAddr_11[32] ?
	       wci_lastConfigAddr_11[31:0] :
	       32'hFFFFFFFF ;
  assign x_data__h105393 = { wci_wReset_n_12, 26'd0, wci_wTimeout_12 } ;
  assign x_data__h105399 =
	     wci_lastConfigAddr_12[32] ?
	       wci_lastConfigAddr_12[31:0] :
	       32'hFFFFFFFF ;
  assign x_data__h105446 = { wci_wReset_n_13, 26'd0, wci_wTimeout_13 } ;
  assign x_data__h105452 =
	     wci_lastConfigAddr_13[32] ?
	       wci_lastConfigAddr_13[31:0] :
	       32'hFFFFFFFF ;
  assign x_data__h105499 = { wci_wReset_n_14, 26'd0, wci_wTimeout_14 } ;
  assign x_data__h105505 =
	     wci_lastConfigAddr_14[32] ?
	       wci_lastConfigAddr_14[31:0] :
	       32'hFFFFFFFF ;
`ifdef not
  assign x_f__h4848 = { timeServ_setRefF$dD_OUT[31:0], 16'h0 } ;
`endif
  always@(wrkAct or
	  wci_respF_14$D_OUT or
	  wci_respF$D_OUT or
	  wci_respF_1$D_OUT or
	  wci_respF_2$D_OUT or
	  wci_respF_3$D_OUT or
	  wci_respF_4$D_OUT or
	  wci_respF_5$D_OUT or
	  wci_respF_6$D_OUT or
	  wci_respF_7$D_OUT or
	  wci_respF_8$D_OUT or
	  wci_respF_9$D_OUT or
	  wci_respF_10$D_OUT or
	  wci_respF_11$D_OUT or wci_respF_12$D_OUT or wci_respF_13$D_OUT)
  begin
    case (wrkAct)
      4'd0: rtnData__h113334 = wci_respF$D_OUT[31:0];
      4'd1: rtnData__h113334 = wci_respF_1$D_OUT[31:0];
      4'd2: rtnData__h113334 = wci_respF_2$D_OUT[31:0];
      4'd3: rtnData__h113334 = wci_respF_3$D_OUT[31:0];
      4'd4: rtnData__h113334 = wci_respF_4$D_OUT[31:0];
      4'd5: rtnData__h113334 = wci_respF_5$D_OUT[31:0];
      4'd6: rtnData__h113334 = wci_respF_6$D_OUT[31:0];
      4'd7: rtnData__h113334 = wci_respF_7$D_OUT[31:0];
      4'd8: rtnData__h113334 = wci_respF_8$D_OUT[31:0];
      4'd9: rtnData__h113334 = wci_respF_9$D_OUT[31:0];
      4'd10: rtnData__h113334 = wci_respF_10$D_OUT[31:0];
      4'd11: rtnData__h113334 = wci_respF_11$D_OUT[31:0];
      4'd12: rtnData__h113334 = wci_respF_12$D_OUT[31:0];
      4'd13: rtnData__h113334 = wci_respF_13$D_OUT[31:0];
      default: rtnData__h113334 = wci_respF_14$D_OUT[31:0];
    endcase
  end
  always@(wrkAct or
	  wci_respF_14$EMPTY_N or
	  wci_respF$EMPTY_N or
	  wci_respF_1$EMPTY_N or
	  wci_respF_2$EMPTY_N or
	  wci_respF_3$EMPTY_N or
	  wci_respF_4$EMPTY_N or
	  wci_respF_5$EMPTY_N or
	  wci_respF_6$EMPTY_N or
	  wci_respF_7$EMPTY_N or
	  wci_respF_8$EMPTY_N or
	  wci_respF_9$EMPTY_N or
	  wci_respF_10$EMPTY_N or
	  wci_respF_11$EMPTY_N or
	  wci_respF_12$EMPTY_N or wci_respF_13$EMPTY_N)
  begin
    case (wrkAct)
      4'd0:
	  IF_wrkAct_077_EQ_0_078_THEN_wci_respF_i_notEmp_ETC___d6132 =
	      wci_respF$EMPTY_N;
      4'd1:
	  IF_wrkAct_077_EQ_0_078_THEN_wci_respF_i_notEmp_ETC___d6132 =
	      wci_respF_1$EMPTY_N;
      4'd2:
	  IF_wrkAct_077_EQ_0_078_THEN_wci_respF_i_notEmp_ETC___d6132 =
	      wci_respF_2$EMPTY_N;
      4'd3:
	  IF_wrkAct_077_EQ_0_078_THEN_wci_respF_i_notEmp_ETC___d6132 =
	      wci_respF_3$EMPTY_N;
      4'd4:
	  IF_wrkAct_077_EQ_0_078_THEN_wci_respF_i_notEmp_ETC___d6132 =
	      wci_respF_4$EMPTY_N;
      4'd5:
	  IF_wrkAct_077_EQ_0_078_THEN_wci_respF_i_notEmp_ETC___d6132 =
	      wci_respF_5$EMPTY_N;
      4'd6:
	  IF_wrkAct_077_EQ_0_078_THEN_wci_respF_i_notEmp_ETC___d6132 =
	      wci_respF_6$EMPTY_N;
      4'd7:
	  IF_wrkAct_077_EQ_0_078_THEN_wci_respF_i_notEmp_ETC___d6132 =
	      wci_respF_7$EMPTY_N;
      4'd8:
	  IF_wrkAct_077_EQ_0_078_THEN_wci_respF_i_notEmp_ETC___d6132 =
	      wci_respF_8$EMPTY_N;
      4'd9:
	  IF_wrkAct_077_EQ_0_078_THEN_wci_respF_i_notEmp_ETC___d6132 =
	      wci_respF_9$EMPTY_N;
      4'd10:
	  IF_wrkAct_077_EQ_0_078_THEN_wci_respF_i_notEmp_ETC___d6132 =
	      wci_respF_10$EMPTY_N;
      4'd11:
	  IF_wrkAct_077_EQ_0_078_THEN_wci_respF_i_notEmp_ETC___d6132 =
	      wci_respF_11$EMPTY_N;
      4'd12:
	  IF_wrkAct_077_EQ_0_078_THEN_wci_respF_i_notEmp_ETC___d6132 =
	      wci_respF_12$EMPTY_N;
      4'd13:
	  IF_wrkAct_077_EQ_0_078_THEN_wci_respF_i_notEmp_ETC___d6132 =
	      wci_respF_13$EMPTY_N;
      default: IF_wrkAct_077_EQ_0_078_THEN_wci_respF_i_notEmp_ETC___d6132 =
		   wrkAct != 4'd14 || wci_respF_14$EMPTY_N;
    endcase
  end
  always@(cpReq or
	  x__h106341 or
`ifdef not
	  pciDevice or
`endif
	  x__h106890 or
	  cpStatus__h75932 or scratch20 or scratch24 or cpControl)
  begin
    case (cpReq[11:4])
      8'h0:
	  IF_cpReq_363_BITS_11_TO_4_366_EQ_0x0_445_THEN__ETC___d6178 =
	      32'h4F70656E;
      8'h04:
	  IF_cpReq_363_BITS_11_TO_4_366_EQ_0x0_445_THEN__ETC___d6178 =
	      32'h43504900;
      8'h08:
	  IF_cpReq_363_BITS_11_TO_4_366_EQ_0x0_445_THEN__ETC___d6178 =
	      32'h00000001;
      8'h0C:
	  IF_cpReq_363_BITS_11_TO_4_366_EQ_0x0_445_THEN__ETC___d6178 =
	      32'd1347452376;
      8'h10:
	  IF_cpReq_363_BITS_11_TO_4_366_EQ_0x0_445_THEN__ETC___d6178 =
	      { 17'd0, x__h106341 };
      8'h14:
	  IF_cpReq_363_BITS_11_TO_4_366_EQ_0x0_445_THEN__ETC___d6178 =
`ifdef not
	      { 16'd0, pciDevice };
`else
	      { 16'd0, 16'd0 };
`endif
      8'h18:
	  IF_cpReq_363_BITS_11_TO_4_366_EQ_0x0_445_THEN__ETC___d6178 =
	      { 17'd0, x__h106890 };
      8'h1C:
	  IF_cpReq_363_BITS_11_TO_4_366_EQ_0x0_445_THEN__ETC___d6178 =
	      cpStatus__h75932;
      8'h20:
	  IF_cpReq_363_BITS_11_TO_4_366_EQ_0x0_445_THEN__ETC___d6178 =
	      scratch20;
      8'h24:
	  IF_cpReq_363_BITS_11_TO_4_366_EQ_0x0_445_THEN__ETC___d6178 =
	      scratch24;
      8'h28:
	  IF_cpReq_363_BITS_11_TO_4_366_EQ_0x0_445_THEN__ETC___d6178 =
	      cpControl;
      default: IF_cpReq_363_BITS_11_TO_4_366_EQ_0x0_445_THEN__ETC___d6178 =
		   32'd0;
    endcase
  end
`ifdef not
  always@(cpReq or
	  timeServ_ppsLostSticky or
	  timeServ_gpsInSticky or
	  timeServ_ppsInSticky or
	  timeServ_timeSetSticky or
	  timeServ_ppsOKCC$dD_OUT or
	  timeServ_ppsLostCC$dD_OUT or
	  timeServ_rollingPPSIn$dD_OUT or
	  timeServ_rplTimeControl or
	  timeServ_nowInCC$dD_OUT or
	  deltaTime or
	  timeServ_refPerPPS$dD_OUT or readCntReg or devDNAV$wget)
  begin
    case (cpReq[11:4])
      8'h30:
	  IF_cpReq_363_BITS_11_TO_4_366_EQ_0x30_595_THEN_ETC___d6177 =
	      { timeServ_ppsLostSticky,
		timeServ_gpsInSticky,
		timeServ_ppsInSticky,
		timeServ_timeSetSticky,
		timeServ_ppsOKCC$dD_OUT,
		timeServ_ppsLostCC$dD_OUT,
		18'h0,
		timeServ_rollingPPSIn$dD_OUT };
      8'h34:
	  IF_cpReq_363_BITS_11_TO_4_366_EQ_0x30_595_THEN_ETC___d6177 =
	      { 27'd0, timeServ_rplTimeControl };
      8'h38:
	  IF_cpReq_363_BITS_11_TO_4_366_EQ_0x30_595_THEN_ETC___d6177 =
	      timeServ_nowInCC$dD_OUT[63:32];
      8'h3C:
	  IF_cpReq_363_BITS_11_TO_4_366_EQ_0x30_595_THEN_ETC___d6177 =
	      timeServ_nowInCC$dD_OUT[31:0];
      8'h40:
	  IF_cpReq_363_BITS_11_TO_4_366_EQ_0x30_595_THEN_ETC___d6177 =
	      deltaTime[63:32];
      8'h44:
	  IF_cpReq_363_BITS_11_TO_4_366_EQ_0x30_595_THEN_ETC___d6177 =
	      deltaTime[31:0];
      8'h48:
	  IF_cpReq_363_BITS_11_TO_4_366_EQ_0x30_595_THEN_ETC___d6177 =
	      { 4'd0, timeServ_refPerPPS$dD_OUT };
      8'h4C:
	  IF_cpReq_363_BITS_11_TO_4_366_EQ_0x30_595_THEN_ETC___d6177 =
	      readCntReg;
      8'h50:
	  IF_cpReq_363_BITS_11_TO_4_366_EQ_0x30_595_THEN_ETC___d6177 =
	      devDNAV$wget[31:0];
      8'h54:
	  IF_cpReq_363_BITS_11_TO_4_366_EQ_0x30_595_THEN_ETC___d6177 =
	      devDNAV$wget[63:32];
      8'h7C:
	  IF_cpReq_363_BITS_11_TO_4_366_EQ_0x30_595_THEN_ETC___d6177 = 32'd2;
      8'h80:
	  IF_cpReq_363_BITS_11_TO_4_366_EQ_0x30_595_THEN_ETC___d6177 =
	      32'd268435464;
      default: IF_cpReq_363_BITS_11_TO_4_366_EQ_0x30_595_THEN_ETC___d6177 =
		   32'd268566536;
    endcase
  end
  always@(cpReq or uuid_arg)
  begin
    case (cpReq[9:6])
      4'd0:
	  CASE_cpReq_BITS_9_TO_6_uuid_arg_BITS_31_TO_0_0_ETC__q3 =
	      uuid_arg[511:480];
      4'd1:
	  CASE_cpReq_BITS_9_TO_6_uuid_arg_BITS_31_TO_0_0_ETC__q3 =
	      uuid_arg[479:448];
      4'd2:
	  CASE_cpReq_BITS_9_TO_6_uuid_arg_BITS_31_TO_0_0_ETC__q3 =
	      uuid_arg[447:416];
      4'd3:
	  CASE_cpReq_BITS_9_TO_6_uuid_arg_BITS_31_TO_0_0_ETC__q3 =
	      uuid_arg[415:384];
      4'd4:
	  CASE_cpReq_BITS_9_TO_6_uuid_arg_BITS_31_TO_0_0_ETC__q3 =
	      uuid_arg[383:352];
      4'd5:
	  CASE_cpReq_BITS_9_TO_6_uuid_arg_BITS_31_TO_0_0_ETC__q3 =
	      uuid_arg[351:320];
      4'd6:
	  CASE_cpReq_BITS_9_TO_6_uuid_arg_BITS_31_TO_0_0_ETC__q3 =
	      uuid_arg[319:288];
      4'd7:
	  CASE_cpReq_BITS_9_TO_6_uuid_arg_BITS_31_TO_0_0_ETC__q3 =
	      uuid_arg[287:256];
      4'h8:
	  CASE_cpReq_BITS_9_TO_6_uuid_arg_BITS_31_TO_0_0_ETC__q3 =
	      uuid_arg[255:224];
      4'h9:
	  CASE_cpReq_BITS_9_TO_6_uuid_arg_BITS_31_TO_0_0_ETC__q3 =
	      uuid_arg[223:192];
      4'hA:
	  CASE_cpReq_BITS_9_TO_6_uuid_arg_BITS_31_TO_0_0_ETC__q3 =
	      uuid_arg[191:160];
      4'd11:
	  CASE_cpReq_BITS_9_TO_6_uuid_arg_BITS_31_TO_0_0_ETC__q3 =
	      uuid_arg[159:128];
      4'hC:
	  CASE_cpReq_BITS_9_TO_6_uuid_arg_BITS_31_TO_0_0_ETC__q3 =
	      uuid_arg[127:96];
      4'd13:
	  CASE_cpReq_BITS_9_TO_6_uuid_arg_BITS_31_TO_0_0_ETC__q3 =
	      uuid_arg[95:64];
      4'd14:
	  CASE_cpReq_BITS_9_TO_6_uuid_arg_BITS_31_TO_0_0_ETC__q3 =
	      uuid_arg[63:32];
      4'd15:
	  CASE_cpReq_BITS_9_TO_6_uuid_arg_BITS_31_TO_0_0_ETC__q3 =
	      uuid_arg[31:0];
    endcase
  end
`endif

  // handling of inlined registers

  always@(posedge CLK)
  begin
    if (RST_N == `BSV_RESET_VALUE)
      begin
        cpControl <= `BSV_ASSIGNMENT_DELAY 32'd0;
	cpReq <= `BSV_ASSIGNMENT_DELAY 65'h02AAAAAAAAAAAAAAA;
`ifdef not
	deltaTime <= `BSV_ASSIGNMENT_DELAY 64'd0;
`endif
	dispatched <= `BSV_ASSIGNMENT_DELAY 1'd0;
`ifdef not
	dna_cnt <= `BSV_ASSIGNMENT_DELAY 7'd0;
	dna_rdReg <= `BSV_ASSIGNMENT_DELAY 1'd0;
	dna_shftReg <= `BSV_ASSIGNMENT_DELAY 1'd0;
	dna_sr <= `BSV_ASSIGNMENT_DELAY 57'd0;
`endif
	readCntReg <= `BSV_ASSIGNMENT_DELAY 32'd0;
	rogueTLP <= `BSV_ASSIGNMENT_DELAY 4'd0;
`ifdef not
	rom_serverAdapter_cnt <= `BSV_ASSIGNMENT_DELAY 3'd0;
	rom_serverAdapter_s1 <= `BSV_ASSIGNMENT_DELAY 2'd0;
`endif
	scratch20 <= `BSV_ASSIGNMENT_DELAY 32'd0;
	scratch24 <= `BSV_ASSIGNMENT_DELAY 32'd0;
`ifdef not
	timeServ_gpsInSticky <= `BSV_ASSIGNMENT_DELAY 1'd0;
	timeServ_ppsInSticky <= `BSV_ASSIGNMENT_DELAY 1'd0;
	timeServ_ppsLostSticky <= `BSV_ASSIGNMENT_DELAY 1'd0;
	timeServ_rplTimeControl <= `BSV_ASSIGNMENT_DELAY 5'd0;
	timeServ_timeSetSticky <= `BSV_ASSIGNMENT_DELAY 1'd0;
`endif
	warmResetP <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_busy <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_busy_1 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_busy_10 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_busy_11 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_busy_12 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_busy_13 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_busy_14 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_busy_2 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_busy_3 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_busy_4 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_busy_5 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_busy_6 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_busy_7 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_busy_8 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_busy_9 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_lastConfigAddr <= `BSV_ASSIGNMENT_DELAY 33'h0AAAAAAAA;
	wci_lastConfigAddr_1 <= `BSV_ASSIGNMENT_DELAY 33'h0AAAAAAAA;
	wci_lastConfigAddr_10 <= `BSV_ASSIGNMENT_DELAY 33'h0AAAAAAAA;
	wci_lastConfigAddr_11 <= `BSV_ASSIGNMENT_DELAY 33'h0AAAAAAAA;
	wci_lastConfigAddr_12 <= `BSV_ASSIGNMENT_DELAY 33'h0AAAAAAAA;
	wci_lastConfigAddr_13 <= `BSV_ASSIGNMENT_DELAY 33'h0AAAAAAAA;
	wci_lastConfigAddr_14 <= `BSV_ASSIGNMENT_DELAY 33'h0AAAAAAAA;
	wci_lastConfigAddr_2 <= `BSV_ASSIGNMENT_DELAY 33'h0AAAAAAAA;
	wci_lastConfigAddr_3 <= `BSV_ASSIGNMENT_DELAY 33'h0AAAAAAAA;
	wci_lastConfigAddr_4 <= `BSV_ASSIGNMENT_DELAY 33'h0AAAAAAAA;
	wci_lastConfigAddr_5 <= `BSV_ASSIGNMENT_DELAY 33'h0AAAAAAAA;
	wci_lastConfigAddr_6 <= `BSV_ASSIGNMENT_DELAY 33'h0AAAAAAAA;
	wci_lastConfigAddr_7 <= `BSV_ASSIGNMENT_DELAY 33'h0AAAAAAAA;
	wci_lastConfigAddr_8 <= `BSV_ASSIGNMENT_DELAY 33'h0AAAAAAAA;
	wci_lastConfigAddr_9 <= `BSV_ASSIGNMENT_DELAY 33'h0AAAAAAAA;
	wci_lastConfigBE <= `BSV_ASSIGNMENT_DELAY 5'd10;
	wci_lastConfigBE_1 <= `BSV_ASSIGNMENT_DELAY 5'd10;
	wci_lastConfigBE_10 <= `BSV_ASSIGNMENT_DELAY 5'd10;
	wci_lastConfigBE_11 <= `BSV_ASSIGNMENT_DELAY 5'd10;
	wci_lastConfigBE_12 <= `BSV_ASSIGNMENT_DELAY 5'd10;
	wci_lastConfigBE_13 <= `BSV_ASSIGNMENT_DELAY 5'd10;
	wci_lastConfigBE_14 <= `BSV_ASSIGNMENT_DELAY 5'd10;
	wci_lastConfigBE_2 <= `BSV_ASSIGNMENT_DELAY 5'd10;
	wci_lastConfigBE_3 <= `BSV_ASSIGNMENT_DELAY 5'd10;
	wci_lastConfigBE_4 <= `BSV_ASSIGNMENT_DELAY 5'd10;
	wci_lastConfigBE_5 <= `BSV_ASSIGNMENT_DELAY 5'd10;
	wci_lastConfigBE_6 <= `BSV_ASSIGNMENT_DELAY 5'd10;
	wci_lastConfigBE_7 <= `BSV_ASSIGNMENT_DELAY 5'd10;
	wci_lastConfigBE_8 <= `BSV_ASSIGNMENT_DELAY 5'd10;
	wci_lastConfigBE_9 <= `BSV_ASSIGNMENT_DELAY 5'd10;
	wci_lastControlOp <= `BSV_ASSIGNMENT_DELAY 4'd2;
	wci_lastControlOp_1 <= `BSV_ASSIGNMENT_DELAY 4'd2;
	wci_lastControlOp_10 <= `BSV_ASSIGNMENT_DELAY 4'd2;
	wci_lastControlOp_11 <= `BSV_ASSIGNMENT_DELAY 4'd2;
	wci_lastControlOp_12 <= `BSV_ASSIGNMENT_DELAY 4'd2;
	wci_lastControlOp_13 <= `BSV_ASSIGNMENT_DELAY 4'd2;
	wci_lastControlOp_14 <= `BSV_ASSIGNMENT_DELAY 4'd2;
	wci_lastControlOp_2 <= `BSV_ASSIGNMENT_DELAY 4'd2;
	wci_lastControlOp_3 <= `BSV_ASSIGNMENT_DELAY 4'd2;
	wci_lastControlOp_4 <= `BSV_ASSIGNMENT_DELAY 4'd2;
	wci_lastControlOp_5 <= `BSV_ASSIGNMENT_DELAY 4'd2;
	wci_lastControlOp_6 <= `BSV_ASSIGNMENT_DELAY 4'd2;
	wci_lastControlOp_7 <= `BSV_ASSIGNMENT_DELAY 4'd2;
	wci_lastControlOp_8 <= `BSV_ASSIGNMENT_DELAY 4'd2;
	wci_lastControlOp_9 <= `BSV_ASSIGNMENT_DELAY 4'd2;
	wci_lastOpWrite <= `BSV_ASSIGNMENT_DELAY 2'd0;
	wci_lastOpWrite_1 <= `BSV_ASSIGNMENT_DELAY 2'd0;
	wci_lastOpWrite_10 <= `BSV_ASSIGNMENT_DELAY 2'd0;
	wci_lastOpWrite_11 <= `BSV_ASSIGNMENT_DELAY 2'd0;
	wci_lastOpWrite_12 <= `BSV_ASSIGNMENT_DELAY 2'd0;
	wci_lastOpWrite_13 <= `BSV_ASSIGNMENT_DELAY 2'd0;
	wci_lastOpWrite_14 <= `BSV_ASSIGNMENT_DELAY 2'd0;
	wci_lastOpWrite_2 <= `BSV_ASSIGNMENT_DELAY 2'd0;
	wci_lastOpWrite_3 <= `BSV_ASSIGNMENT_DELAY 2'd0;
	wci_lastOpWrite_4 <= `BSV_ASSIGNMENT_DELAY 2'd0;
	wci_lastOpWrite_5 <= `BSV_ASSIGNMENT_DELAY 2'd0;
	wci_lastOpWrite_6 <= `BSV_ASSIGNMENT_DELAY 2'd0;
	wci_lastOpWrite_7 <= `BSV_ASSIGNMENT_DELAY 2'd0;
	wci_lastOpWrite_8 <= `BSV_ASSIGNMENT_DELAY 2'd0;
	wci_lastOpWrite_9 <= `BSV_ASSIGNMENT_DELAY 2'd0;
	wci_mFlagReg <= `BSV_ASSIGNMENT_DELAY 2'b10;
	wci_mFlagReg_1 <= `BSV_ASSIGNMENT_DELAY 2'b10;
	wci_mFlagReg_10 <= `BSV_ASSIGNMENT_DELAY 2'b10;
	wci_mFlagReg_11 <= `BSV_ASSIGNMENT_DELAY 2'b10;
	wci_mFlagReg_12 <= `BSV_ASSIGNMENT_DELAY 2'b10;
	wci_mFlagReg_13 <= `BSV_ASSIGNMENT_DELAY 2'b10;
	wci_mFlagReg_14 <= `BSV_ASSIGNMENT_DELAY 2'b10;
	wci_mFlagReg_2 <= `BSV_ASSIGNMENT_DELAY 2'b10;
	wci_mFlagReg_3 <= `BSV_ASSIGNMENT_DELAY 2'b10;
	wci_mFlagReg_4 <= `BSV_ASSIGNMENT_DELAY 2'b10;
	wci_mFlagReg_5 <= `BSV_ASSIGNMENT_DELAY 2'b10;
	wci_mFlagReg_6 <= `BSV_ASSIGNMENT_DELAY 2'b10;
	wci_mFlagReg_7 <= `BSV_ASSIGNMENT_DELAY 2'b10;
	wci_mFlagReg_8 <= `BSV_ASSIGNMENT_DELAY 2'b10;
	wci_mFlagReg_9 <= `BSV_ASSIGNMENT_DELAY 2'b10;
	wci_pageWindow <= `BSV_ASSIGNMENT_DELAY 12'd0;
	wci_pageWindow_1 <= `BSV_ASSIGNMENT_DELAY 12'd0;
	wci_pageWindow_10 <= `BSV_ASSIGNMENT_DELAY 12'd0;
	wci_pageWindow_11 <= `BSV_ASSIGNMENT_DELAY 12'd0;
	wci_pageWindow_12 <= `BSV_ASSIGNMENT_DELAY 12'd0;
	wci_pageWindow_13 <= `BSV_ASSIGNMENT_DELAY 12'd0;
	wci_pageWindow_14 <= `BSV_ASSIGNMENT_DELAY 12'd0;
	wci_pageWindow_2 <= `BSV_ASSIGNMENT_DELAY 12'd0;
	wci_pageWindow_3 <= `BSV_ASSIGNMENT_DELAY 12'd0;
	wci_pageWindow_4 <= `BSV_ASSIGNMENT_DELAY 12'd0;
	wci_pageWindow_5 <= `BSV_ASSIGNMENT_DELAY 12'd0;
	wci_pageWindow_6 <= `BSV_ASSIGNMENT_DELAY 12'd0;
	wci_pageWindow_7 <= `BSV_ASSIGNMENT_DELAY 12'd0;
	wci_pageWindow_8 <= `BSV_ASSIGNMENT_DELAY 12'd0;
	wci_pageWindow_9 <= `BSV_ASSIGNMENT_DELAY 12'd0;
	wci_reqERR <= `BSV_ASSIGNMENT_DELAY 3'd0;
	wci_reqERR_1 <= `BSV_ASSIGNMENT_DELAY 3'd0;
	wci_reqERR_10 <= `BSV_ASSIGNMENT_DELAY 3'd0;
	wci_reqERR_11 <= `BSV_ASSIGNMENT_DELAY 3'd0;
	wci_reqERR_12 <= `BSV_ASSIGNMENT_DELAY 3'd0;
	wci_reqERR_13 <= `BSV_ASSIGNMENT_DELAY 3'd0;
	wci_reqERR_14 <= `BSV_ASSIGNMENT_DELAY 3'd0;
	wci_reqERR_2 <= `BSV_ASSIGNMENT_DELAY 3'd0;
	wci_reqERR_3 <= `BSV_ASSIGNMENT_DELAY 3'd0;
	wci_reqERR_4 <= `BSV_ASSIGNMENT_DELAY 3'd0;
	wci_reqERR_5 <= `BSV_ASSIGNMENT_DELAY 3'd0;
	wci_reqERR_6 <= `BSV_ASSIGNMENT_DELAY 3'd0;
	wci_reqERR_7 <= `BSV_ASSIGNMENT_DELAY 3'd0;
	wci_reqERR_8 <= `BSV_ASSIGNMENT_DELAY 3'd0;
	wci_reqERR_9 <= `BSV_ASSIGNMENT_DELAY 3'd0;
	wci_reqFAIL <= `BSV_ASSIGNMENT_DELAY 3'd0;
	wci_reqFAIL_1 <= `BSV_ASSIGNMENT_DELAY 3'd0;
	wci_reqFAIL_10 <= `BSV_ASSIGNMENT_DELAY 3'd0;
	wci_reqFAIL_11 <= `BSV_ASSIGNMENT_DELAY 3'd0;
	wci_reqFAIL_12 <= `BSV_ASSIGNMENT_DELAY 3'd0;
	wci_reqFAIL_13 <= `BSV_ASSIGNMENT_DELAY 3'd0;
	wci_reqFAIL_14 <= `BSV_ASSIGNMENT_DELAY 3'd0;
	wci_reqFAIL_2 <= `BSV_ASSIGNMENT_DELAY 3'd0;
	wci_reqFAIL_3 <= `BSV_ASSIGNMENT_DELAY 3'd0;
	wci_reqFAIL_4 <= `BSV_ASSIGNMENT_DELAY 3'd0;
	wci_reqFAIL_5 <= `BSV_ASSIGNMENT_DELAY 3'd0;
	wci_reqFAIL_6 <= `BSV_ASSIGNMENT_DELAY 3'd0;
	wci_reqFAIL_7 <= `BSV_ASSIGNMENT_DELAY 3'd0;
	wci_reqFAIL_8 <= `BSV_ASSIGNMENT_DELAY 3'd0;
	wci_reqFAIL_9 <= `BSV_ASSIGNMENT_DELAY 3'd0;
	wci_reqF_10_c_r <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_reqF_10_q_0 <= `BSV_ASSIGNMENT_DELAY 72'h0000000000AAAAAAAA;
	wci_reqF_11_c_r <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_reqF_11_q_0 <= `BSV_ASSIGNMENT_DELAY 72'h0000000000AAAAAAAA;
	wci_reqF_12_c_r <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_reqF_12_q_0 <= `BSV_ASSIGNMENT_DELAY 72'h0000000000AAAAAAAA;
	wci_reqF_13_c_r <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_reqF_13_q_0 <= `BSV_ASSIGNMENT_DELAY 72'h0000000000AAAAAAAA;
	wci_reqF_14_c_r <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_reqF_14_q_0 <= `BSV_ASSIGNMENT_DELAY 72'h0000000000AAAAAAAA;
	wci_reqF_1_c_r <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_reqF_1_q_0 <= `BSV_ASSIGNMENT_DELAY 72'h0000000000AAAAAAAA;
	wci_reqF_2_c_r <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_reqF_2_q_0 <= `BSV_ASSIGNMENT_DELAY 72'h0000000000AAAAAAAA;
	wci_reqF_3_c_r <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_reqF_3_q_0 <= `BSV_ASSIGNMENT_DELAY 72'h0000000000AAAAAAAA;
	wci_reqF_4_c_r <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_reqF_4_q_0 <= `BSV_ASSIGNMENT_DELAY 72'h0000000000AAAAAAAA;
	wci_reqF_5_c_r <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_reqF_5_q_0 <= `BSV_ASSIGNMENT_DELAY 72'h0000000000AAAAAAAA;
	wci_reqF_6_c_r <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_reqF_6_q_0 <= `BSV_ASSIGNMENT_DELAY 72'h0000000000AAAAAAAA;
	wci_reqF_7_c_r <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_reqF_7_q_0 <= `BSV_ASSIGNMENT_DELAY 72'h0000000000AAAAAAAA;
	wci_reqF_8_c_r <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_reqF_8_q_0 <= `BSV_ASSIGNMENT_DELAY 72'h0000000000AAAAAAAA;
	wci_reqF_9_c_r <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_reqF_9_q_0 <= `BSV_ASSIGNMENT_DELAY 72'h0000000000AAAAAAAA;
	wci_reqF_c_r <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_reqF_q_0 <= `BSV_ASSIGNMENT_DELAY 72'h0000000000AAAAAAAA;
	wci_reqPend <= `BSV_ASSIGNMENT_DELAY 2'd0;
	wci_reqPend_1 <= `BSV_ASSIGNMENT_DELAY 2'd0;
	wci_reqPend_10 <= `BSV_ASSIGNMENT_DELAY 2'd0;
	wci_reqPend_11 <= `BSV_ASSIGNMENT_DELAY 2'd0;
	wci_reqPend_12 <= `BSV_ASSIGNMENT_DELAY 2'd0;
	wci_reqPend_13 <= `BSV_ASSIGNMENT_DELAY 2'd0;
	wci_reqPend_14 <= `BSV_ASSIGNMENT_DELAY 2'd0;
	wci_reqPend_2 <= `BSV_ASSIGNMENT_DELAY 2'd0;
	wci_reqPend_3 <= `BSV_ASSIGNMENT_DELAY 2'd0;
	wci_reqPend_4 <= `BSV_ASSIGNMENT_DELAY 2'd0;
	wci_reqPend_5 <= `BSV_ASSIGNMENT_DELAY 2'd0;
	wci_reqPend_6 <= `BSV_ASSIGNMENT_DELAY 2'd0;
	wci_reqPend_7 <= `BSV_ASSIGNMENT_DELAY 2'd0;
	wci_reqPend_8 <= `BSV_ASSIGNMENT_DELAY 2'd0;
	wci_reqPend_9 <= `BSV_ASSIGNMENT_DELAY 2'd0;
	wci_reqTO <= `BSV_ASSIGNMENT_DELAY 3'd0;
	wci_reqTO_1 <= `BSV_ASSIGNMENT_DELAY 3'd0;
	wci_reqTO_10 <= `BSV_ASSIGNMENT_DELAY 3'd0;
	wci_reqTO_11 <= `BSV_ASSIGNMENT_DELAY 3'd0;
	wci_reqTO_12 <= `BSV_ASSIGNMENT_DELAY 3'd0;
	wci_reqTO_13 <= `BSV_ASSIGNMENT_DELAY 3'd0;
	wci_reqTO_14 <= `BSV_ASSIGNMENT_DELAY 3'd0;
	wci_reqTO_2 <= `BSV_ASSIGNMENT_DELAY 3'd0;
	wci_reqTO_3 <= `BSV_ASSIGNMENT_DELAY 3'd0;
	wci_reqTO_4 <= `BSV_ASSIGNMENT_DELAY 3'd0;
	wci_reqTO_5 <= `BSV_ASSIGNMENT_DELAY 3'd0;
	wci_reqTO_6 <= `BSV_ASSIGNMENT_DELAY 3'd0;
	wci_reqTO_7 <= `BSV_ASSIGNMENT_DELAY 3'd0;
	wci_reqTO_8 <= `BSV_ASSIGNMENT_DELAY 3'd0;
	wci_reqTO_9 <= `BSV_ASSIGNMENT_DELAY 3'd0;
	wci_respTimr <= `BSV_ASSIGNMENT_DELAY 32'd0;
	wci_respTimrAct <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_respTimrAct_1 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_respTimrAct_10 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_respTimrAct_11 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_respTimrAct_12 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_respTimrAct_13 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_respTimrAct_14 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_respTimrAct_2 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_respTimrAct_3 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_respTimrAct_4 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_respTimrAct_5 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_respTimrAct_6 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_respTimrAct_7 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_respTimrAct_8 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_respTimrAct_9 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_respTimr_1 <= `BSV_ASSIGNMENT_DELAY 32'd0;
	wci_respTimr_10 <= `BSV_ASSIGNMENT_DELAY 32'd0;
	wci_respTimr_11 <= `BSV_ASSIGNMENT_DELAY 32'd0;
	wci_respTimr_12 <= `BSV_ASSIGNMENT_DELAY 32'd0;
	wci_respTimr_13 <= `BSV_ASSIGNMENT_DELAY 32'd0;
	wci_respTimr_14 <= `BSV_ASSIGNMENT_DELAY 32'd0;
	wci_respTimr_2 <= `BSV_ASSIGNMENT_DELAY 32'd0;
	wci_respTimr_3 <= `BSV_ASSIGNMENT_DELAY 32'd0;
	wci_respTimr_4 <= `BSV_ASSIGNMENT_DELAY 32'd0;
	wci_respTimr_5 <= `BSV_ASSIGNMENT_DELAY 32'd0;
	wci_respTimr_6 <= `BSV_ASSIGNMENT_DELAY 32'd0;
	wci_respTimr_7 <= `BSV_ASSIGNMENT_DELAY 32'd0;
	wci_respTimr_8 <= `BSV_ASSIGNMENT_DELAY 32'd0;
	wci_respTimr_9 <= `BSV_ASSIGNMENT_DELAY 32'd0;
	wci_sThreadBusy_d <= `BSV_ASSIGNMENT_DELAY 1'd1;
	wci_sThreadBusy_d_1 <= `BSV_ASSIGNMENT_DELAY 1'd1;
	wci_sThreadBusy_d_10 <= `BSV_ASSIGNMENT_DELAY 1'd1;
	wci_sThreadBusy_d_11 <= `BSV_ASSIGNMENT_DELAY 1'd1;
	wci_sThreadBusy_d_12 <= `BSV_ASSIGNMENT_DELAY 1'd1;
	wci_sThreadBusy_d_13 <= `BSV_ASSIGNMENT_DELAY 1'd1;
	wci_sThreadBusy_d_14 <= `BSV_ASSIGNMENT_DELAY 1'd1;
	wci_sThreadBusy_d_2 <= `BSV_ASSIGNMENT_DELAY 1'd1;
	wci_sThreadBusy_d_3 <= `BSV_ASSIGNMENT_DELAY 1'd1;
	wci_sThreadBusy_d_4 <= `BSV_ASSIGNMENT_DELAY 1'd1;
	wci_sThreadBusy_d_5 <= `BSV_ASSIGNMENT_DELAY 1'd1;
	wci_sThreadBusy_d_6 <= `BSV_ASSIGNMENT_DELAY 1'd1;
	wci_sThreadBusy_d_7 <= `BSV_ASSIGNMENT_DELAY 1'd1;
	wci_sThreadBusy_d_8 <= `BSV_ASSIGNMENT_DELAY 1'd1;
	wci_sThreadBusy_d_9 <= `BSV_ASSIGNMENT_DELAY 1'd1;
	wci_sfCap <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_sfCapClear <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_sfCapClear_10 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_sfCapClear_11 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_sfCapClear_12 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_sfCapClear_13 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_sfCapClear_14 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_sfCapClear_1_1 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_sfCapClear_2 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_sfCapClear_3 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_sfCapClear_4 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_sfCapClear_5 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_sfCapClear_6 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_sfCapClear_7 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_sfCapClear_8 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_sfCapClear_9 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_sfCapSet <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_sfCapSet_10 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_sfCapSet_11 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_sfCapSet_12 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_sfCapSet_13 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_sfCapSet_14 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_sfCapSet_1_1 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_sfCapSet_2 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_sfCapSet_3 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_sfCapSet_4 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_sfCapSet_5 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_sfCapSet_6 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_sfCapSet_7 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_sfCapSet_8 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_sfCapSet_9 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_sfCap_1 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_sfCap_10 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_sfCap_11 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_sfCap_12 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_sfCap_13 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_sfCap_14 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_sfCap_2 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_sfCap_3 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_sfCap_4 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_sfCap_5 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_sfCap_6 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_sfCap_7 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_sfCap_8 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_sfCap_9 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_slvPresent <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_slvPresent_1 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_slvPresent_10 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_slvPresent_11 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_slvPresent_12 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_slvPresent_13 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_slvPresent_14 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_slvPresent_2 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_slvPresent_3 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_slvPresent_4 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_slvPresent_5 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_slvPresent_6 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_slvPresent_7 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_slvPresent_8 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_slvPresent_9 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_wReset_n <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_wReset_n_1 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_wReset_n_10 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_wReset_n_11 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_wReset_n_12 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_wReset_n_13 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_wReset_n_14 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_wReset_n_2 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_wReset_n_3 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_wReset_n_4 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_wReset_n_5 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_wReset_n_6 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_wReset_n_7 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_wReset_n_8 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_wReset_n_9 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wci_wTimeout <= `BSV_ASSIGNMENT_DELAY 5'h04;
	wci_wTimeout_1 <= `BSV_ASSIGNMENT_DELAY 5'h04;
	wci_wTimeout_10 <= `BSV_ASSIGNMENT_DELAY 5'h04;
	wci_wTimeout_11 <= `BSV_ASSIGNMENT_DELAY 5'h04;
	wci_wTimeout_12 <= `BSV_ASSIGNMENT_DELAY 5'h04;
	wci_wTimeout_13 <= `BSV_ASSIGNMENT_DELAY 5'h04;
	wci_wTimeout_14 <= `BSV_ASSIGNMENT_DELAY 5'h04;
	wci_wTimeout_2 <= `BSV_ASSIGNMENT_DELAY 5'h04;
	wci_wTimeout_3 <= `BSV_ASSIGNMENT_DELAY 5'h04;
	wci_wTimeout_4 <= `BSV_ASSIGNMENT_DELAY 5'h04;
	wci_wTimeout_5 <= `BSV_ASSIGNMENT_DELAY 5'h04;
	wci_wTimeout_6 <= `BSV_ASSIGNMENT_DELAY 5'h04;
	wci_wTimeout_7 <= `BSV_ASSIGNMENT_DELAY 5'h04;
	wci_wTimeout_8 <= `BSV_ASSIGNMENT_DELAY 5'h04;
	wci_wTimeout_9 <= `BSV_ASSIGNMENT_DELAY 5'h04;
	wrkAct <= `BSV_ASSIGNMENT_DELAY 4'd0;
      end
    else
      begin
        if (cpControl$EN) cpControl <= `BSV_ASSIGNMENT_DELAY cpControl$D_IN;
	if (cpReq$EN) cpReq <= `BSV_ASSIGNMENT_DELAY cpReq$D_IN;
`ifdef not
	if (deltaTime$EN) deltaTime <= `BSV_ASSIGNMENT_DELAY deltaTime$D_IN;
`endif
	if (dispatched$EN)
	  dispatched <= `BSV_ASSIGNMENT_DELAY dispatched$D_IN;
`ifdef not
	if (dna_cnt$EN) dna_cnt <= `BSV_ASSIGNMENT_DELAY dna_cnt$D_IN;
	if (dna_rdReg$EN) dna_rdReg <= `BSV_ASSIGNMENT_DELAY dna_rdReg$D_IN;
	if (dna_shftReg$EN)
	  dna_shftReg <= `BSV_ASSIGNMENT_DELAY dna_shftReg$D_IN;
	if (dna_sr$EN) dna_sr <= `BSV_ASSIGNMENT_DELAY dna_sr$D_IN;
`endif
	if (readCntReg$EN)
	  readCntReg <= `BSV_ASSIGNMENT_DELAY readCntReg$D_IN;
	if (rogueTLP$EN) rogueTLP <= `BSV_ASSIGNMENT_DELAY rogueTLP$D_IN;
`ifdef not
	if (rom_serverAdapter_cnt$EN)
	  rom_serverAdapter_cnt <= `BSV_ASSIGNMENT_DELAY
	      rom_serverAdapter_cnt$D_IN;
	if (rom_serverAdapter_s1$EN)
	  rom_serverAdapter_s1 <= `BSV_ASSIGNMENT_DELAY
	      rom_serverAdapter_s1$D_IN;
`endif
	if (scratch20$EN) scratch20 <= `BSV_ASSIGNMENT_DELAY scratch20$D_IN;
	if (scratch24$EN) scratch24 <= `BSV_ASSIGNMENT_DELAY scratch24$D_IN;
`ifdef not
	if (timeServ_gpsInSticky$EN)
	  timeServ_gpsInSticky <= `BSV_ASSIGNMENT_DELAY
	      timeServ_gpsInSticky$D_IN;
	if (timeServ_ppsInSticky$EN)
	  timeServ_ppsInSticky <= `BSV_ASSIGNMENT_DELAY
	      timeServ_ppsInSticky$D_IN;
	if (timeServ_ppsLostSticky$EN)
	  timeServ_ppsLostSticky <= `BSV_ASSIGNMENT_DELAY
	      timeServ_ppsLostSticky$D_IN;
	if (timeServ_rplTimeControl$EN)
	  timeServ_rplTimeControl <= `BSV_ASSIGNMENT_DELAY
	      timeServ_rplTimeControl$D_IN;
	if (timeServ_timeSetSticky$EN)
	  timeServ_timeSetSticky <= `BSV_ASSIGNMENT_DELAY
	      timeServ_timeSetSticky$D_IN;
`endif
	if (warmResetP$EN)
	  warmResetP <= `BSV_ASSIGNMENT_DELAY warmResetP$D_IN;
	if (wci_busy$EN) wci_busy <= `BSV_ASSIGNMENT_DELAY wci_busy$D_IN;
	if (wci_busy_1$EN)
	  wci_busy_1 <= `BSV_ASSIGNMENT_DELAY wci_busy_1$D_IN;
	if (wci_busy_10$EN)
	  wci_busy_10 <= `BSV_ASSIGNMENT_DELAY wci_busy_10$D_IN;
	if (wci_busy_11$EN)
	  wci_busy_11 <= `BSV_ASSIGNMENT_DELAY wci_busy_11$D_IN;
	if (wci_busy_12$EN)
	  wci_busy_12 <= `BSV_ASSIGNMENT_DELAY wci_busy_12$D_IN;
	if (wci_busy_13$EN)
	  wci_busy_13 <= `BSV_ASSIGNMENT_DELAY wci_busy_13$D_IN;
	if (wci_busy_14$EN)
	  wci_busy_14 <= `BSV_ASSIGNMENT_DELAY wci_busy_14$D_IN;
	if (wci_busy_2$EN)
	  wci_busy_2 <= `BSV_ASSIGNMENT_DELAY wci_busy_2$D_IN;
	if (wci_busy_3$EN)
	  wci_busy_3 <= `BSV_ASSIGNMENT_DELAY wci_busy_3$D_IN;
	if (wci_busy_4$EN)
	  wci_busy_4 <= `BSV_ASSIGNMENT_DELAY wci_busy_4$D_IN;
	if (wci_busy_5$EN)
	  wci_busy_5 <= `BSV_ASSIGNMENT_DELAY wci_busy_5$D_IN;
	if (wci_busy_6$EN)
	  wci_busy_6 <= `BSV_ASSIGNMENT_DELAY wci_busy_6$D_IN;
	if (wci_busy_7$EN)
	  wci_busy_7 <= `BSV_ASSIGNMENT_DELAY wci_busy_7$D_IN;
	if (wci_busy_8$EN)
	  wci_busy_8 <= `BSV_ASSIGNMENT_DELAY wci_busy_8$D_IN;
	if (wci_busy_9$EN)
	  wci_busy_9 <= `BSV_ASSIGNMENT_DELAY wci_busy_9$D_IN;
	if (wci_lastConfigAddr$EN)
	  wci_lastConfigAddr <= `BSV_ASSIGNMENT_DELAY wci_lastConfigAddr$D_IN;
	if (wci_lastConfigAddr_1$EN)
	  wci_lastConfigAddr_1 <= `BSV_ASSIGNMENT_DELAY
	      wci_lastConfigAddr_1$D_IN;
	if (wci_lastConfigAddr_10$EN)
	  wci_lastConfigAddr_10 <= `BSV_ASSIGNMENT_DELAY
	      wci_lastConfigAddr_10$D_IN;
	if (wci_lastConfigAddr_11$EN)
	  wci_lastConfigAddr_11 <= `BSV_ASSIGNMENT_DELAY
	      wci_lastConfigAddr_11$D_IN;
	if (wci_lastConfigAddr_12$EN)
	  wci_lastConfigAddr_12 <= `BSV_ASSIGNMENT_DELAY
	      wci_lastConfigAddr_12$D_IN;
	if (wci_lastConfigAddr_13$EN)
	  wci_lastConfigAddr_13 <= `BSV_ASSIGNMENT_DELAY
	      wci_lastConfigAddr_13$D_IN;
	if (wci_lastConfigAddr_14$EN)
	  wci_lastConfigAddr_14 <= `BSV_ASSIGNMENT_DELAY
	      wci_lastConfigAddr_14$D_IN;
	if (wci_lastConfigAddr_2$EN)
	  wci_lastConfigAddr_2 <= `BSV_ASSIGNMENT_DELAY
	      wci_lastConfigAddr_2$D_IN;
	if (wci_lastConfigAddr_3$EN)
	  wci_lastConfigAddr_3 <= `BSV_ASSIGNMENT_DELAY
	      wci_lastConfigAddr_3$D_IN;
	if (wci_lastConfigAddr_4$EN)
	  wci_lastConfigAddr_4 <= `BSV_ASSIGNMENT_DELAY
	      wci_lastConfigAddr_4$D_IN;
	if (wci_lastConfigAddr_5$EN)
	  wci_lastConfigAddr_5 <= `BSV_ASSIGNMENT_DELAY
	      wci_lastConfigAddr_5$D_IN;
	if (wci_lastConfigAddr_6$EN)
	  wci_lastConfigAddr_6 <= `BSV_ASSIGNMENT_DELAY
	      wci_lastConfigAddr_6$D_IN;
	if (wci_lastConfigAddr_7$EN)
	  wci_lastConfigAddr_7 <= `BSV_ASSIGNMENT_DELAY
	      wci_lastConfigAddr_7$D_IN;
	if (wci_lastConfigAddr_8$EN)
	  wci_lastConfigAddr_8 <= `BSV_ASSIGNMENT_DELAY
	      wci_lastConfigAddr_8$D_IN;
	if (wci_lastConfigAddr_9$EN)
	  wci_lastConfigAddr_9 <= `BSV_ASSIGNMENT_DELAY
	      wci_lastConfigAddr_9$D_IN;
	if (wci_lastConfigBE$EN)
	  wci_lastConfigBE <= `BSV_ASSIGNMENT_DELAY wci_lastConfigBE$D_IN;
	if (wci_lastConfigBE_1$EN)
	  wci_lastConfigBE_1 <= `BSV_ASSIGNMENT_DELAY wci_lastConfigBE_1$D_IN;
	if (wci_lastConfigBE_10$EN)
	  wci_lastConfigBE_10 <= `BSV_ASSIGNMENT_DELAY
	      wci_lastConfigBE_10$D_IN;
	if (wci_lastConfigBE_11$EN)
	  wci_lastConfigBE_11 <= `BSV_ASSIGNMENT_DELAY
	      wci_lastConfigBE_11$D_IN;
	if (wci_lastConfigBE_12$EN)
	  wci_lastConfigBE_12 <= `BSV_ASSIGNMENT_DELAY
	      wci_lastConfigBE_12$D_IN;
	if (wci_lastConfigBE_13$EN)
	  wci_lastConfigBE_13 <= `BSV_ASSIGNMENT_DELAY
	      wci_lastConfigBE_13$D_IN;
	if (wci_lastConfigBE_14$EN)
	  wci_lastConfigBE_14 <= `BSV_ASSIGNMENT_DELAY
	      wci_lastConfigBE_14$D_IN;
	if (wci_lastConfigBE_2$EN)
	  wci_lastConfigBE_2 <= `BSV_ASSIGNMENT_DELAY wci_lastConfigBE_2$D_IN;
	if (wci_lastConfigBE_3$EN)
	  wci_lastConfigBE_3 <= `BSV_ASSIGNMENT_DELAY wci_lastConfigBE_3$D_IN;
	if (wci_lastConfigBE_4$EN)
	  wci_lastConfigBE_4 <= `BSV_ASSIGNMENT_DELAY wci_lastConfigBE_4$D_IN;
	if (wci_lastConfigBE_5$EN)
	  wci_lastConfigBE_5 <= `BSV_ASSIGNMENT_DELAY wci_lastConfigBE_5$D_IN;
	if (wci_lastConfigBE_6$EN)
	  wci_lastConfigBE_6 <= `BSV_ASSIGNMENT_DELAY wci_lastConfigBE_6$D_IN;
	if (wci_lastConfigBE_7$EN)
	  wci_lastConfigBE_7 <= `BSV_ASSIGNMENT_DELAY wci_lastConfigBE_7$D_IN;
	if (wci_lastConfigBE_8$EN)
	  wci_lastConfigBE_8 <= `BSV_ASSIGNMENT_DELAY wci_lastConfigBE_8$D_IN;
	if (wci_lastConfigBE_9$EN)
	  wci_lastConfigBE_9 <= `BSV_ASSIGNMENT_DELAY wci_lastConfigBE_9$D_IN;
	if (wci_lastControlOp$EN)
	  wci_lastControlOp <= `BSV_ASSIGNMENT_DELAY wci_lastControlOp$D_IN;
	if (wci_lastControlOp_1$EN)
	  wci_lastControlOp_1 <= `BSV_ASSIGNMENT_DELAY
	      wci_lastControlOp_1$D_IN;
	if (wci_lastControlOp_10$EN)
	  wci_lastControlOp_10 <= `BSV_ASSIGNMENT_DELAY
	      wci_lastControlOp_10$D_IN;
	if (wci_lastControlOp_11$EN)
	  wci_lastControlOp_11 <= `BSV_ASSIGNMENT_DELAY
	      wci_lastControlOp_11$D_IN;
	if (wci_lastControlOp_12$EN)
	  wci_lastControlOp_12 <= `BSV_ASSIGNMENT_DELAY
	      wci_lastControlOp_12$D_IN;
	if (wci_lastControlOp_13$EN)
	  wci_lastControlOp_13 <= `BSV_ASSIGNMENT_DELAY
	      wci_lastControlOp_13$D_IN;
	if (wci_lastControlOp_14$EN)
	  wci_lastControlOp_14 <= `BSV_ASSIGNMENT_DELAY
	      wci_lastControlOp_14$D_IN;
	if (wci_lastControlOp_2$EN)
	  wci_lastControlOp_2 <= `BSV_ASSIGNMENT_DELAY
	      wci_lastControlOp_2$D_IN;
	if (wci_lastControlOp_3$EN)
	  wci_lastControlOp_3 <= `BSV_ASSIGNMENT_DELAY
	      wci_lastControlOp_3$D_IN;
	if (wci_lastControlOp_4$EN)
	  wci_lastControlOp_4 <= `BSV_ASSIGNMENT_DELAY
	      wci_lastControlOp_4$D_IN;
	if (wci_lastControlOp_5$EN)
	  wci_lastControlOp_5 <= `BSV_ASSIGNMENT_DELAY
	      wci_lastControlOp_5$D_IN;
	if (wci_lastControlOp_6$EN)
	  wci_lastControlOp_6 <= `BSV_ASSIGNMENT_DELAY
	      wci_lastControlOp_6$D_IN;
	if (wci_lastControlOp_7$EN)
	  wci_lastControlOp_7 <= `BSV_ASSIGNMENT_DELAY
	      wci_lastControlOp_7$D_IN;
	if (wci_lastControlOp_8$EN)
	  wci_lastControlOp_8 <= `BSV_ASSIGNMENT_DELAY
	      wci_lastControlOp_8$D_IN;
	if (wci_lastControlOp_9$EN)
	  wci_lastControlOp_9 <= `BSV_ASSIGNMENT_DELAY
	      wci_lastControlOp_9$D_IN;
	if (wci_lastOpWrite$EN)
	  wci_lastOpWrite <= `BSV_ASSIGNMENT_DELAY wci_lastOpWrite$D_IN;
	if (wci_lastOpWrite_1$EN)
	  wci_lastOpWrite_1 <= `BSV_ASSIGNMENT_DELAY wci_lastOpWrite_1$D_IN;
	if (wci_lastOpWrite_10$EN)
	  wci_lastOpWrite_10 <= `BSV_ASSIGNMENT_DELAY wci_lastOpWrite_10$D_IN;
	if (wci_lastOpWrite_11$EN)
	  wci_lastOpWrite_11 <= `BSV_ASSIGNMENT_DELAY wci_lastOpWrite_11$D_IN;
	if (wci_lastOpWrite_12$EN)
	  wci_lastOpWrite_12 <= `BSV_ASSIGNMENT_DELAY wci_lastOpWrite_12$D_IN;
	if (wci_lastOpWrite_13$EN)
	  wci_lastOpWrite_13 <= `BSV_ASSIGNMENT_DELAY wci_lastOpWrite_13$D_IN;
	if (wci_lastOpWrite_14$EN)
	  wci_lastOpWrite_14 <= `BSV_ASSIGNMENT_DELAY wci_lastOpWrite_14$D_IN;
	if (wci_lastOpWrite_2$EN)
	  wci_lastOpWrite_2 <= `BSV_ASSIGNMENT_DELAY wci_lastOpWrite_2$D_IN;
	if (wci_lastOpWrite_3$EN)
	  wci_lastOpWrite_3 <= `BSV_ASSIGNMENT_DELAY wci_lastOpWrite_3$D_IN;
	if (wci_lastOpWrite_4$EN)
	  wci_lastOpWrite_4 <= `BSV_ASSIGNMENT_DELAY wci_lastOpWrite_4$D_IN;
	if (wci_lastOpWrite_5$EN)
	  wci_lastOpWrite_5 <= `BSV_ASSIGNMENT_DELAY wci_lastOpWrite_5$D_IN;
	if (wci_lastOpWrite_6$EN)
	  wci_lastOpWrite_6 <= `BSV_ASSIGNMENT_DELAY wci_lastOpWrite_6$D_IN;
	if (wci_lastOpWrite_7$EN)
	  wci_lastOpWrite_7 <= `BSV_ASSIGNMENT_DELAY wci_lastOpWrite_7$D_IN;
	if (wci_lastOpWrite_8$EN)
	  wci_lastOpWrite_8 <= `BSV_ASSIGNMENT_DELAY wci_lastOpWrite_8$D_IN;
	if (wci_lastOpWrite_9$EN)
	  wci_lastOpWrite_9 <= `BSV_ASSIGNMENT_DELAY wci_lastOpWrite_9$D_IN;
	if (wci_mFlagReg$EN)
	  wci_mFlagReg <= `BSV_ASSIGNMENT_DELAY wci_mFlagReg$D_IN;
	if (wci_mFlagReg_1$EN)
	  wci_mFlagReg_1 <= `BSV_ASSIGNMENT_DELAY wci_mFlagReg_1$D_IN;
	if (wci_mFlagReg_10$EN)
	  wci_mFlagReg_10 <= `BSV_ASSIGNMENT_DELAY wci_mFlagReg_10$D_IN;
	if (wci_mFlagReg_11$EN)
	  wci_mFlagReg_11 <= `BSV_ASSIGNMENT_DELAY wci_mFlagReg_11$D_IN;
	if (wci_mFlagReg_12$EN)
	  wci_mFlagReg_12 <= `BSV_ASSIGNMENT_DELAY wci_mFlagReg_12$D_IN;
	if (wci_mFlagReg_13$EN)
	  wci_mFlagReg_13 <= `BSV_ASSIGNMENT_DELAY wci_mFlagReg_13$D_IN;
	if (wci_mFlagReg_14$EN)
	  wci_mFlagReg_14 <= `BSV_ASSIGNMENT_DELAY wci_mFlagReg_14$D_IN;
	if (wci_mFlagReg_2$EN)
	  wci_mFlagReg_2 <= `BSV_ASSIGNMENT_DELAY wci_mFlagReg_2$D_IN;
	if (wci_mFlagReg_3$EN)
	  wci_mFlagReg_3 <= `BSV_ASSIGNMENT_DELAY wci_mFlagReg_3$D_IN;
	if (wci_mFlagReg_4$EN)
	  wci_mFlagReg_4 <= `BSV_ASSIGNMENT_DELAY wci_mFlagReg_4$D_IN;
	if (wci_mFlagReg_5$EN)
	  wci_mFlagReg_5 <= `BSV_ASSIGNMENT_DELAY wci_mFlagReg_5$D_IN;
	if (wci_mFlagReg_6$EN)
	  wci_mFlagReg_6 <= `BSV_ASSIGNMENT_DELAY wci_mFlagReg_6$D_IN;
	if (wci_mFlagReg_7$EN)
	  wci_mFlagReg_7 <= `BSV_ASSIGNMENT_DELAY wci_mFlagReg_7$D_IN;
	if (wci_mFlagReg_8$EN)
	  wci_mFlagReg_8 <= `BSV_ASSIGNMENT_DELAY wci_mFlagReg_8$D_IN;
	if (wci_mFlagReg_9$EN)
	  wci_mFlagReg_9 <= `BSV_ASSIGNMENT_DELAY wci_mFlagReg_9$D_IN;
	if (wci_pageWindow$EN)
	  wci_pageWindow <= `BSV_ASSIGNMENT_DELAY wci_pageWindow$D_IN;
	if (wci_pageWindow_1$EN)
	  wci_pageWindow_1 <= `BSV_ASSIGNMENT_DELAY wci_pageWindow_1$D_IN;
	if (wci_pageWindow_10$EN)
	  wci_pageWindow_10 <= `BSV_ASSIGNMENT_DELAY wci_pageWindow_10$D_IN;
	if (wci_pageWindow_11$EN)
	  wci_pageWindow_11 <= `BSV_ASSIGNMENT_DELAY wci_pageWindow_11$D_IN;
	if (wci_pageWindow_12$EN)
	  wci_pageWindow_12 <= `BSV_ASSIGNMENT_DELAY wci_pageWindow_12$D_IN;
	if (wci_pageWindow_13$EN)
	  wci_pageWindow_13 <= `BSV_ASSIGNMENT_DELAY wci_pageWindow_13$D_IN;
	if (wci_pageWindow_14$EN)
	  wci_pageWindow_14 <= `BSV_ASSIGNMENT_DELAY wci_pageWindow_14$D_IN;
	if (wci_pageWindow_2$EN)
	  wci_pageWindow_2 <= `BSV_ASSIGNMENT_DELAY wci_pageWindow_2$D_IN;
	if (wci_pageWindow_3$EN)
	  wci_pageWindow_3 <= `BSV_ASSIGNMENT_DELAY wci_pageWindow_3$D_IN;
	if (wci_pageWindow_4$EN)
	  wci_pageWindow_4 <= `BSV_ASSIGNMENT_DELAY wci_pageWindow_4$D_IN;
	if (wci_pageWindow_5$EN)
	  wci_pageWindow_5 <= `BSV_ASSIGNMENT_DELAY wci_pageWindow_5$D_IN;
	if (wci_pageWindow_6$EN)
	  wci_pageWindow_6 <= `BSV_ASSIGNMENT_DELAY wci_pageWindow_6$D_IN;
	if (wci_pageWindow_7$EN)
	  wci_pageWindow_7 <= `BSV_ASSIGNMENT_DELAY wci_pageWindow_7$D_IN;
	if (wci_pageWindow_8$EN)
	  wci_pageWindow_8 <= `BSV_ASSIGNMENT_DELAY wci_pageWindow_8$D_IN;
	if (wci_pageWindow_9$EN)
	  wci_pageWindow_9 <= `BSV_ASSIGNMENT_DELAY wci_pageWindow_9$D_IN;
	if (wci_reqERR$EN)
	  wci_reqERR <= `BSV_ASSIGNMENT_DELAY wci_reqERR$D_IN;
	if (wci_reqERR_1$EN)
	  wci_reqERR_1 <= `BSV_ASSIGNMENT_DELAY wci_reqERR_1$D_IN;
	if (wci_reqERR_10$EN)
	  wci_reqERR_10 <= `BSV_ASSIGNMENT_DELAY wci_reqERR_10$D_IN;
	if (wci_reqERR_11$EN)
	  wci_reqERR_11 <= `BSV_ASSIGNMENT_DELAY wci_reqERR_11$D_IN;
	if (wci_reqERR_12$EN)
	  wci_reqERR_12 <= `BSV_ASSIGNMENT_DELAY wci_reqERR_12$D_IN;
	if (wci_reqERR_13$EN)
	  wci_reqERR_13 <= `BSV_ASSIGNMENT_DELAY wci_reqERR_13$D_IN;
	if (wci_reqERR_14$EN)
	  wci_reqERR_14 <= `BSV_ASSIGNMENT_DELAY wci_reqERR_14$D_IN;
	if (wci_reqERR_2$EN)
	  wci_reqERR_2 <= `BSV_ASSIGNMENT_DELAY wci_reqERR_2$D_IN;
	if (wci_reqERR_3$EN)
	  wci_reqERR_3 <= `BSV_ASSIGNMENT_DELAY wci_reqERR_3$D_IN;
	if (wci_reqERR_4$EN)
	  wci_reqERR_4 <= `BSV_ASSIGNMENT_DELAY wci_reqERR_4$D_IN;
	if (wci_reqERR_5$EN)
	  wci_reqERR_5 <= `BSV_ASSIGNMENT_DELAY wci_reqERR_5$D_IN;
	if (wci_reqERR_6$EN)
	  wci_reqERR_6 <= `BSV_ASSIGNMENT_DELAY wci_reqERR_6$D_IN;
	if (wci_reqERR_7$EN)
	  wci_reqERR_7 <= `BSV_ASSIGNMENT_DELAY wci_reqERR_7$D_IN;
	if (wci_reqERR_8$EN)
	  wci_reqERR_8 <= `BSV_ASSIGNMENT_DELAY wci_reqERR_8$D_IN;
	if (wci_reqERR_9$EN)
	  wci_reqERR_9 <= `BSV_ASSIGNMENT_DELAY wci_reqERR_9$D_IN;
	if (wci_reqFAIL$EN)
	  wci_reqFAIL <= `BSV_ASSIGNMENT_DELAY wci_reqFAIL$D_IN;
	if (wci_reqFAIL_1$EN)
	  wci_reqFAIL_1 <= `BSV_ASSIGNMENT_DELAY wci_reqFAIL_1$D_IN;
	if (wci_reqFAIL_10$EN)
	  wci_reqFAIL_10 <= `BSV_ASSIGNMENT_DELAY wci_reqFAIL_10$D_IN;
	if (wci_reqFAIL_11$EN)
	  wci_reqFAIL_11 <= `BSV_ASSIGNMENT_DELAY wci_reqFAIL_11$D_IN;
	if (wci_reqFAIL_12$EN)
	  wci_reqFAIL_12 <= `BSV_ASSIGNMENT_DELAY wci_reqFAIL_12$D_IN;
	if (wci_reqFAIL_13$EN)
	  wci_reqFAIL_13 <= `BSV_ASSIGNMENT_DELAY wci_reqFAIL_13$D_IN;
	if (wci_reqFAIL_14$EN)
	  wci_reqFAIL_14 <= `BSV_ASSIGNMENT_DELAY wci_reqFAIL_14$D_IN;
	if (wci_reqFAIL_2$EN)
	  wci_reqFAIL_2 <= `BSV_ASSIGNMENT_DELAY wci_reqFAIL_2$D_IN;
	if (wci_reqFAIL_3$EN)
	  wci_reqFAIL_3 <= `BSV_ASSIGNMENT_DELAY wci_reqFAIL_3$D_IN;
	if (wci_reqFAIL_4$EN)
	  wci_reqFAIL_4 <= `BSV_ASSIGNMENT_DELAY wci_reqFAIL_4$D_IN;
	if (wci_reqFAIL_5$EN)
	  wci_reqFAIL_5 <= `BSV_ASSIGNMENT_DELAY wci_reqFAIL_5$D_IN;
	if (wci_reqFAIL_6$EN)
	  wci_reqFAIL_6 <= `BSV_ASSIGNMENT_DELAY wci_reqFAIL_6$D_IN;
	if (wci_reqFAIL_7$EN)
	  wci_reqFAIL_7 <= `BSV_ASSIGNMENT_DELAY wci_reqFAIL_7$D_IN;
	if (wci_reqFAIL_8$EN)
	  wci_reqFAIL_8 <= `BSV_ASSIGNMENT_DELAY wci_reqFAIL_8$D_IN;
	if (wci_reqFAIL_9$EN)
	  wci_reqFAIL_9 <= `BSV_ASSIGNMENT_DELAY wci_reqFAIL_9$D_IN;
	if (wci_reqF_10_c_r$EN)
	  wci_reqF_10_c_r <= `BSV_ASSIGNMENT_DELAY wci_reqF_10_c_r$D_IN;
	if (wci_reqF_10_q_0$EN)
	  wci_reqF_10_q_0 <= `BSV_ASSIGNMENT_DELAY wci_reqF_10_q_0$D_IN;
	if (wci_reqF_11_c_r$EN)
	  wci_reqF_11_c_r <= `BSV_ASSIGNMENT_DELAY wci_reqF_11_c_r$D_IN;
	if (wci_reqF_11_q_0$EN)
	  wci_reqF_11_q_0 <= `BSV_ASSIGNMENT_DELAY wci_reqF_11_q_0$D_IN;
	if (wci_reqF_12_c_r$EN)
	  wci_reqF_12_c_r <= `BSV_ASSIGNMENT_DELAY wci_reqF_12_c_r$D_IN;
	if (wci_reqF_12_q_0$EN)
	  wci_reqF_12_q_0 <= `BSV_ASSIGNMENT_DELAY wci_reqF_12_q_0$D_IN;
	if (wci_reqF_13_c_r$EN)
	  wci_reqF_13_c_r <= `BSV_ASSIGNMENT_DELAY wci_reqF_13_c_r$D_IN;
	if (wci_reqF_13_q_0$EN)
	  wci_reqF_13_q_0 <= `BSV_ASSIGNMENT_DELAY wci_reqF_13_q_0$D_IN;
	if (wci_reqF_14_c_r$EN)
	  wci_reqF_14_c_r <= `BSV_ASSIGNMENT_DELAY wci_reqF_14_c_r$D_IN;
	if (wci_reqF_14_q_0$EN)
	  wci_reqF_14_q_0 <= `BSV_ASSIGNMENT_DELAY wci_reqF_14_q_0$D_IN;
	if (wci_reqF_1_c_r$EN)
	  wci_reqF_1_c_r <= `BSV_ASSIGNMENT_DELAY wci_reqF_1_c_r$D_IN;
	if (wci_reqF_1_q_0$EN)
	  wci_reqF_1_q_0 <= `BSV_ASSIGNMENT_DELAY wci_reqF_1_q_0$D_IN;
	if (wci_reqF_2_c_r$EN)
	  wci_reqF_2_c_r <= `BSV_ASSIGNMENT_DELAY wci_reqF_2_c_r$D_IN;
	if (wci_reqF_2_q_0$EN)
	  wci_reqF_2_q_0 <= `BSV_ASSIGNMENT_DELAY wci_reqF_2_q_0$D_IN;
	if (wci_reqF_3_c_r$EN)
	  wci_reqF_3_c_r <= `BSV_ASSIGNMENT_DELAY wci_reqF_3_c_r$D_IN;
	if (wci_reqF_3_q_0$EN)
	  wci_reqF_3_q_0 <= `BSV_ASSIGNMENT_DELAY wci_reqF_3_q_0$D_IN;
	if (wci_reqF_4_c_r$EN)
	  wci_reqF_4_c_r <= `BSV_ASSIGNMENT_DELAY wci_reqF_4_c_r$D_IN;
	if (wci_reqF_4_q_0$EN)
	  wci_reqF_4_q_0 <= `BSV_ASSIGNMENT_DELAY wci_reqF_4_q_0$D_IN;
	if (wci_reqF_5_c_r$EN)
	  wci_reqF_5_c_r <= `BSV_ASSIGNMENT_DELAY wci_reqF_5_c_r$D_IN;
	if (wci_reqF_5_q_0$EN)
	  wci_reqF_5_q_0 <= `BSV_ASSIGNMENT_DELAY wci_reqF_5_q_0$D_IN;
	if (wci_reqF_6_c_r$EN)
	  wci_reqF_6_c_r <= `BSV_ASSIGNMENT_DELAY wci_reqF_6_c_r$D_IN;
	if (wci_reqF_6_q_0$EN)
	  wci_reqF_6_q_0 <= `BSV_ASSIGNMENT_DELAY wci_reqF_6_q_0$D_IN;
	if (wci_reqF_7_c_r$EN)
	  wci_reqF_7_c_r <= `BSV_ASSIGNMENT_DELAY wci_reqF_7_c_r$D_IN;
	if (wci_reqF_7_q_0$EN)
	  wci_reqF_7_q_0 <= `BSV_ASSIGNMENT_DELAY wci_reqF_7_q_0$D_IN;
	if (wci_reqF_8_c_r$EN)
	  wci_reqF_8_c_r <= `BSV_ASSIGNMENT_DELAY wci_reqF_8_c_r$D_IN;
	if (wci_reqF_8_q_0$EN)
	  wci_reqF_8_q_0 <= `BSV_ASSIGNMENT_DELAY wci_reqF_8_q_0$D_IN;
	if (wci_reqF_9_c_r$EN)
	  wci_reqF_9_c_r <= `BSV_ASSIGNMENT_DELAY wci_reqF_9_c_r$D_IN;
	if (wci_reqF_9_q_0$EN)
	  wci_reqF_9_q_0 <= `BSV_ASSIGNMENT_DELAY wci_reqF_9_q_0$D_IN;
	if (wci_reqF_c_r$EN)
	  wci_reqF_c_r <= `BSV_ASSIGNMENT_DELAY wci_reqF_c_r$D_IN;
	if (wci_reqF_q_0$EN)
	  wci_reqF_q_0 <= `BSV_ASSIGNMENT_DELAY wci_reqF_q_0$D_IN;
	if (wci_reqPend$EN)
	  wci_reqPend <= `BSV_ASSIGNMENT_DELAY wci_reqPend$D_IN;
	if (wci_reqPend_1$EN)
	  wci_reqPend_1 <= `BSV_ASSIGNMENT_DELAY wci_reqPend_1$D_IN;
	if (wci_reqPend_10$EN)
	  wci_reqPend_10 <= `BSV_ASSIGNMENT_DELAY wci_reqPend_10$D_IN;
	if (wci_reqPend_11$EN)
	  wci_reqPend_11 <= `BSV_ASSIGNMENT_DELAY wci_reqPend_11$D_IN;
	if (wci_reqPend_12$EN)
	  wci_reqPend_12 <= `BSV_ASSIGNMENT_DELAY wci_reqPend_12$D_IN;
	if (wci_reqPend_13$EN)
	  wci_reqPend_13 <= `BSV_ASSIGNMENT_DELAY wci_reqPend_13$D_IN;
	if (wci_reqPend_14$EN)
	  wci_reqPend_14 <= `BSV_ASSIGNMENT_DELAY wci_reqPend_14$D_IN;
	if (wci_reqPend_2$EN)
	  wci_reqPend_2 <= `BSV_ASSIGNMENT_DELAY wci_reqPend_2$D_IN;
	if (wci_reqPend_3$EN)
	  wci_reqPend_3 <= `BSV_ASSIGNMENT_DELAY wci_reqPend_3$D_IN;
	if (wci_reqPend_4$EN)
	  wci_reqPend_4 <= `BSV_ASSIGNMENT_DELAY wci_reqPend_4$D_IN;
	if (wci_reqPend_5$EN)
	  wci_reqPend_5 <= `BSV_ASSIGNMENT_DELAY wci_reqPend_5$D_IN;
	if (wci_reqPend_6$EN)
	  wci_reqPend_6 <= `BSV_ASSIGNMENT_DELAY wci_reqPend_6$D_IN;
	if (wci_reqPend_7$EN)
	  wci_reqPend_7 <= `BSV_ASSIGNMENT_DELAY wci_reqPend_7$D_IN;
	if (wci_reqPend_8$EN)
	  wci_reqPend_8 <= `BSV_ASSIGNMENT_DELAY wci_reqPend_8$D_IN;
	if (wci_reqPend_9$EN)
	  wci_reqPend_9 <= `BSV_ASSIGNMENT_DELAY wci_reqPend_9$D_IN;
	if (wci_reqTO$EN) wci_reqTO <= `BSV_ASSIGNMENT_DELAY wci_reqTO$D_IN;
	if (wci_reqTO_1$EN)
	  wci_reqTO_1 <= `BSV_ASSIGNMENT_DELAY wci_reqTO_1$D_IN;
	if (wci_reqTO_10$EN)
	  wci_reqTO_10 <= `BSV_ASSIGNMENT_DELAY wci_reqTO_10$D_IN;
	if (wci_reqTO_11$EN)
	  wci_reqTO_11 <= `BSV_ASSIGNMENT_DELAY wci_reqTO_11$D_IN;
	if (wci_reqTO_12$EN)
	  wci_reqTO_12 <= `BSV_ASSIGNMENT_DELAY wci_reqTO_12$D_IN;
	if (wci_reqTO_13$EN)
	  wci_reqTO_13 <= `BSV_ASSIGNMENT_DELAY wci_reqTO_13$D_IN;
	if (wci_reqTO_14$EN)
	  wci_reqTO_14 <= `BSV_ASSIGNMENT_DELAY wci_reqTO_14$D_IN;
	if (wci_reqTO_2$EN)
	  wci_reqTO_2 <= `BSV_ASSIGNMENT_DELAY wci_reqTO_2$D_IN;
	if (wci_reqTO_3$EN)
	  wci_reqTO_3 <= `BSV_ASSIGNMENT_DELAY wci_reqTO_3$D_IN;
	if (wci_reqTO_4$EN)
	  wci_reqTO_4 <= `BSV_ASSIGNMENT_DELAY wci_reqTO_4$D_IN;
	if (wci_reqTO_5$EN)
	  wci_reqTO_5 <= `BSV_ASSIGNMENT_DELAY wci_reqTO_5$D_IN;
	if (wci_reqTO_6$EN)
	  wci_reqTO_6 <= `BSV_ASSIGNMENT_DELAY wci_reqTO_6$D_IN;
	if (wci_reqTO_7$EN)
	  wci_reqTO_7 <= `BSV_ASSIGNMENT_DELAY wci_reqTO_7$D_IN;
	if (wci_reqTO_8$EN)
	  wci_reqTO_8 <= `BSV_ASSIGNMENT_DELAY wci_reqTO_8$D_IN;
	if (wci_reqTO_9$EN)
	  wci_reqTO_9 <= `BSV_ASSIGNMENT_DELAY wci_reqTO_9$D_IN;
	if (wci_respTimr$EN)
	  wci_respTimr <= `BSV_ASSIGNMENT_DELAY wci_respTimr$D_IN;
	if (wci_respTimrAct$EN)
	  wci_respTimrAct <= `BSV_ASSIGNMENT_DELAY wci_respTimrAct$D_IN;
	if (wci_respTimrAct_1$EN)
	  wci_respTimrAct_1 <= `BSV_ASSIGNMENT_DELAY wci_respTimrAct_1$D_IN;
	if (wci_respTimrAct_10$EN)
	  wci_respTimrAct_10 <= `BSV_ASSIGNMENT_DELAY wci_respTimrAct_10$D_IN;
	if (wci_respTimrAct_11$EN)
	  wci_respTimrAct_11 <= `BSV_ASSIGNMENT_DELAY wci_respTimrAct_11$D_IN;
	if (wci_respTimrAct_12$EN)
	  wci_respTimrAct_12 <= `BSV_ASSIGNMENT_DELAY wci_respTimrAct_12$D_IN;
	if (wci_respTimrAct_13$EN)
	  wci_respTimrAct_13 <= `BSV_ASSIGNMENT_DELAY wci_respTimrAct_13$D_IN;
	if (wci_respTimrAct_14$EN)
	  wci_respTimrAct_14 <= `BSV_ASSIGNMENT_DELAY wci_respTimrAct_14$D_IN;
	if (wci_respTimrAct_2$EN)
	  wci_respTimrAct_2 <= `BSV_ASSIGNMENT_DELAY wci_respTimrAct_2$D_IN;
	if (wci_respTimrAct_3$EN)
	  wci_respTimrAct_3 <= `BSV_ASSIGNMENT_DELAY wci_respTimrAct_3$D_IN;
	if (wci_respTimrAct_4$EN)
	  wci_respTimrAct_4 <= `BSV_ASSIGNMENT_DELAY wci_respTimrAct_4$D_IN;
	if (wci_respTimrAct_5$EN)
	  wci_respTimrAct_5 <= `BSV_ASSIGNMENT_DELAY wci_respTimrAct_5$D_IN;
	if (wci_respTimrAct_6$EN)
	  wci_respTimrAct_6 <= `BSV_ASSIGNMENT_DELAY wci_respTimrAct_6$D_IN;
	if (wci_respTimrAct_7$EN)
	  wci_respTimrAct_7 <= `BSV_ASSIGNMENT_DELAY wci_respTimrAct_7$D_IN;
	if (wci_respTimrAct_8$EN)
	  wci_respTimrAct_8 <= `BSV_ASSIGNMENT_DELAY wci_respTimrAct_8$D_IN;
	if (wci_respTimrAct_9$EN)
	  wci_respTimrAct_9 <= `BSV_ASSIGNMENT_DELAY wci_respTimrAct_9$D_IN;
	if (wci_respTimr_1$EN)
	  wci_respTimr_1 <= `BSV_ASSIGNMENT_DELAY wci_respTimr_1$D_IN;
	if (wci_respTimr_10$EN)
	  wci_respTimr_10 <= `BSV_ASSIGNMENT_DELAY wci_respTimr_10$D_IN;
	if (wci_respTimr_11$EN)
	  wci_respTimr_11 <= `BSV_ASSIGNMENT_DELAY wci_respTimr_11$D_IN;
	if (wci_respTimr_12$EN)
	  wci_respTimr_12 <= `BSV_ASSIGNMENT_DELAY wci_respTimr_12$D_IN;
	if (wci_respTimr_13$EN)
	  wci_respTimr_13 <= `BSV_ASSIGNMENT_DELAY wci_respTimr_13$D_IN;
	if (wci_respTimr_14$EN)
	  wci_respTimr_14 <= `BSV_ASSIGNMENT_DELAY wci_respTimr_14$D_IN;
	if (wci_respTimr_2$EN)
	  wci_respTimr_2 <= `BSV_ASSIGNMENT_DELAY wci_respTimr_2$D_IN;
	if (wci_respTimr_3$EN)
	  wci_respTimr_3 <= `BSV_ASSIGNMENT_DELAY wci_respTimr_3$D_IN;
	if (wci_respTimr_4$EN)
	  wci_respTimr_4 <= `BSV_ASSIGNMENT_DELAY wci_respTimr_4$D_IN;
	if (wci_respTimr_5$EN)
	  wci_respTimr_5 <= `BSV_ASSIGNMENT_DELAY wci_respTimr_5$D_IN;
	if (wci_respTimr_6$EN)
	  wci_respTimr_6 <= `BSV_ASSIGNMENT_DELAY wci_respTimr_6$D_IN;
	if (wci_respTimr_7$EN)
	  wci_respTimr_7 <= `BSV_ASSIGNMENT_DELAY wci_respTimr_7$D_IN;
	if (wci_respTimr_8$EN)
	  wci_respTimr_8 <= `BSV_ASSIGNMENT_DELAY wci_respTimr_8$D_IN;
	if (wci_respTimr_9$EN)
	  wci_respTimr_9 <= `BSV_ASSIGNMENT_DELAY wci_respTimr_9$D_IN;
	if (wci_sThreadBusy_d$EN)
	  wci_sThreadBusy_d <= `BSV_ASSIGNMENT_DELAY wci_sThreadBusy_d$D_IN;
	if (wci_sThreadBusy_d_1$EN)
	  wci_sThreadBusy_d_1 <= `BSV_ASSIGNMENT_DELAY
	      wci_sThreadBusy_d_1$D_IN;
	if (wci_sThreadBusy_d_10$EN)
	  wci_sThreadBusy_d_10 <= `BSV_ASSIGNMENT_DELAY
	      wci_sThreadBusy_d_10$D_IN;
	if (wci_sThreadBusy_d_11$EN)
	  wci_sThreadBusy_d_11 <= `BSV_ASSIGNMENT_DELAY
	      wci_sThreadBusy_d_11$D_IN;
	if (wci_sThreadBusy_d_12$EN)
	  wci_sThreadBusy_d_12 <= `BSV_ASSIGNMENT_DELAY
	      wci_sThreadBusy_d_12$D_IN;
	if (wci_sThreadBusy_d_13$EN)
	  wci_sThreadBusy_d_13 <= `BSV_ASSIGNMENT_DELAY
	      wci_sThreadBusy_d_13$D_IN;
	if (wci_sThreadBusy_d_14$EN)
	  wci_sThreadBusy_d_14 <= `BSV_ASSIGNMENT_DELAY
	      wci_sThreadBusy_d_14$D_IN;
	if (wci_sThreadBusy_d_2$EN)
	  wci_sThreadBusy_d_2 <= `BSV_ASSIGNMENT_DELAY
	      wci_sThreadBusy_d_2$D_IN;
	if (wci_sThreadBusy_d_3$EN)
	  wci_sThreadBusy_d_3 <= `BSV_ASSIGNMENT_DELAY
	      wci_sThreadBusy_d_3$D_IN;
	if (wci_sThreadBusy_d_4$EN)
	  wci_sThreadBusy_d_4 <= `BSV_ASSIGNMENT_DELAY
	      wci_sThreadBusy_d_4$D_IN;
	if (wci_sThreadBusy_d_5$EN)
	  wci_sThreadBusy_d_5 <= `BSV_ASSIGNMENT_DELAY
	      wci_sThreadBusy_d_5$D_IN;
	if (wci_sThreadBusy_d_6$EN)
	  wci_sThreadBusy_d_6 <= `BSV_ASSIGNMENT_DELAY
	      wci_sThreadBusy_d_6$D_IN;
	if (wci_sThreadBusy_d_7$EN)
	  wci_sThreadBusy_d_7 <= `BSV_ASSIGNMENT_DELAY
	      wci_sThreadBusy_d_7$D_IN;
	if (wci_sThreadBusy_d_8$EN)
	  wci_sThreadBusy_d_8 <= `BSV_ASSIGNMENT_DELAY
	      wci_sThreadBusy_d_8$D_IN;
	if (wci_sThreadBusy_d_9$EN)
	  wci_sThreadBusy_d_9 <= `BSV_ASSIGNMENT_DELAY
	      wci_sThreadBusy_d_9$D_IN;
	if (wci_sfCap$EN) wci_sfCap <= `BSV_ASSIGNMENT_DELAY wci_sfCap$D_IN;
	if (wci_sfCapClear$EN)
	  wci_sfCapClear <= `BSV_ASSIGNMENT_DELAY wci_sfCapClear$D_IN;
	if (wci_sfCapClear_10$EN)
	  wci_sfCapClear_10 <= `BSV_ASSIGNMENT_DELAY wci_sfCapClear_10$D_IN;
	if (wci_sfCapClear_11$EN)
	  wci_sfCapClear_11 <= `BSV_ASSIGNMENT_DELAY wci_sfCapClear_11$D_IN;
	if (wci_sfCapClear_12$EN)
	  wci_sfCapClear_12 <= `BSV_ASSIGNMENT_DELAY wci_sfCapClear_12$D_IN;
	if (wci_sfCapClear_13$EN)
	  wci_sfCapClear_13 <= `BSV_ASSIGNMENT_DELAY wci_sfCapClear_13$D_IN;
	if (wci_sfCapClear_14$EN)
	  wci_sfCapClear_14 <= `BSV_ASSIGNMENT_DELAY wci_sfCapClear_14$D_IN;
	if (wci_sfCapClear_1_1$EN)
	  wci_sfCapClear_1_1 <= `BSV_ASSIGNMENT_DELAY wci_sfCapClear_1_1$D_IN;
	if (wci_sfCapClear_2$EN)
	  wci_sfCapClear_2 <= `BSV_ASSIGNMENT_DELAY wci_sfCapClear_2$D_IN;
	if (wci_sfCapClear_3$EN)
	  wci_sfCapClear_3 <= `BSV_ASSIGNMENT_DELAY wci_sfCapClear_3$D_IN;
	if (wci_sfCapClear_4$EN)
	  wci_sfCapClear_4 <= `BSV_ASSIGNMENT_DELAY wci_sfCapClear_4$D_IN;
	if (wci_sfCapClear_5$EN)
	  wci_sfCapClear_5 <= `BSV_ASSIGNMENT_DELAY wci_sfCapClear_5$D_IN;
	if (wci_sfCapClear_6$EN)
	  wci_sfCapClear_6 <= `BSV_ASSIGNMENT_DELAY wci_sfCapClear_6$D_IN;
	if (wci_sfCapClear_7$EN)
	  wci_sfCapClear_7 <= `BSV_ASSIGNMENT_DELAY wci_sfCapClear_7$D_IN;
	if (wci_sfCapClear_8$EN)
	  wci_sfCapClear_8 <= `BSV_ASSIGNMENT_DELAY wci_sfCapClear_8$D_IN;
	if (wci_sfCapClear_9$EN)
	  wci_sfCapClear_9 <= `BSV_ASSIGNMENT_DELAY wci_sfCapClear_9$D_IN;
	if (wci_sfCapSet$EN)
	  wci_sfCapSet <= `BSV_ASSIGNMENT_DELAY wci_sfCapSet$D_IN;
	if (wci_sfCapSet_10$EN)
	  wci_sfCapSet_10 <= `BSV_ASSIGNMENT_DELAY wci_sfCapSet_10$D_IN;
	if (wci_sfCapSet_11$EN)
	  wci_sfCapSet_11 <= `BSV_ASSIGNMENT_DELAY wci_sfCapSet_11$D_IN;
	if (wci_sfCapSet_12$EN)
	  wci_sfCapSet_12 <= `BSV_ASSIGNMENT_DELAY wci_sfCapSet_12$D_IN;
	if (wci_sfCapSet_13$EN)
	  wci_sfCapSet_13 <= `BSV_ASSIGNMENT_DELAY wci_sfCapSet_13$D_IN;
	if (wci_sfCapSet_14$EN)
	  wci_sfCapSet_14 <= `BSV_ASSIGNMENT_DELAY wci_sfCapSet_14$D_IN;
	if (wci_sfCapSet_1_1$EN)
	  wci_sfCapSet_1_1 <= `BSV_ASSIGNMENT_DELAY wci_sfCapSet_1_1$D_IN;
	if (wci_sfCapSet_2$EN)
	  wci_sfCapSet_2 <= `BSV_ASSIGNMENT_DELAY wci_sfCapSet_2$D_IN;
	if (wci_sfCapSet_3$EN)
	  wci_sfCapSet_3 <= `BSV_ASSIGNMENT_DELAY wci_sfCapSet_3$D_IN;
	if (wci_sfCapSet_4$EN)
	  wci_sfCapSet_4 <= `BSV_ASSIGNMENT_DELAY wci_sfCapSet_4$D_IN;
	if (wci_sfCapSet_5$EN)
	  wci_sfCapSet_5 <= `BSV_ASSIGNMENT_DELAY wci_sfCapSet_5$D_IN;
	if (wci_sfCapSet_6$EN)
	  wci_sfCapSet_6 <= `BSV_ASSIGNMENT_DELAY wci_sfCapSet_6$D_IN;
	if (wci_sfCapSet_7$EN)
	  wci_sfCapSet_7 <= `BSV_ASSIGNMENT_DELAY wci_sfCapSet_7$D_IN;
	if (wci_sfCapSet_8$EN)
	  wci_sfCapSet_8 <= `BSV_ASSIGNMENT_DELAY wci_sfCapSet_8$D_IN;
	if (wci_sfCapSet_9$EN)
	  wci_sfCapSet_9 <= `BSV_ASSIGNMENT_DELAY wci_sfCapSet_9$D_IN;
	if (wci_sfCap_1$EN)
	  wci_sfCap_1 <= `BSV_ASSIGNMENT_DELAY wci_sfCap_1$D_IN;
	if (wci_sfCap_10$EN)
	  wci_sfCap_10 <= `BSV_ASSIGNMENT_DELAY wci_sfCap_10$D_IN;
	if (wci_sfCap_11$EN)
	  wci_sfCap_11 <= `BSV_ASSIGNMENT_DELAY wci_sfCap_11$D_IN;
	if (wci_sfCap_12$EN)
	  wci_sfCap_12 <= `BSV_ASSIGNMENT_DELAY wci_sfCap_12$D_IN;
	if (wci_sfCap_13$EN)
	  wci_sfCap_13 <= `BSV_ASSIGNMENT_DELAY wci_sfCap_13$D_IN;
	if (wci_sfCap_14$EN)
	  wci_sfCap_14 <= `BSV_ASSIGNMENT_DELAY wci_sfCap_14$D_IN;
	if (wci_sfCap_2$EN)
	  wci_sfCap_2 <= `BSV_ASSIGNMENT_DELAY wci_sfCap_2$D_IN;
	if (wci_sfCap_3$EN)
	  wci_sfCap_3 <= `BSV_ASSIGNMENT_DELAY wci_sfCap_3$D_IN;
	if (wci_sfCap_4$EN)
	  wci_sfCap_4 <= `BSV_ASSIGNMENT_DELAY wci_sfCap_4$D_IN;
	if (wci_sfCap_5$EN)
	  wci_sfCap_5 <= `BSV_ASSIGNMENT_DELAY wci_sfCap_5$D_IN;
	if (wci_sfCap_6$EN)
	  wci_sfCap_6 <= `BSV_ASSIGNMENT_DELAY wci_sfCap_6$D_IN;
	if (wci_sfCap_7$EN)
	  wci_sfCap_7 <= `BSV_ASSIGNMENT_DELAY wci_sfCap_7$D_IN;
	if (wci_sfCap_8$EN)
	  wci_sfCap_8 <= `BSV_ASSIGNMENT_DELAY wci_sfCap_8$D_IN;
	if (wci_sfCap_9$EN)
	  wci_sfCap_9 <= `BSV_ASSIGNMENT_DELAY wci_sfCap_9$D_IN;
	if (wci_slvPresent$EN)
	  wci_slvPresent <= `BSV_ASSIGNMENT_DELAY wci_slvPresent$D_IN;
	if (wci_slvPresent_1$EN)
	  wci_slvPresent_1 <= `BSV_ASSIGNMENT_DELAY wci_slvPresent_1$D_IN;
	if (wci_slvPresent_10$EN)
	  wci_slvPresent_10 <= `BSV_ASSIGNMENT_DELAY wci_slvPresent_10$D_IN;
	if (wci_slvPresent_11$EN)
	  wci_slvPresent_11 <= `BSV_ASSIGNMENT_DELAY wci_slvPresent_11$D_IN;
	if (wci_slvPresent_12$EN)
	  wci_slvPresent_12 <= `BSV_ASSIGNMENT_DELAY wci_slvPresent_12$D_IN;
	if (wci_slvPresent_13$EN)
	  wci_slvPresent_13 <= `BSV_ASSIGNMENT_DELAY wci_slvPresent_13$D_IN;
	if (wci_slvPresent_14$EN)
	  wci_slvPresent_14 <= `BSV_ASSIGNMENT_DELAY wci_slvPresent_14$D_IN;
	if (wci_slvPresent_2$EN)
	  wci_slvPresent_2 <= `BSV_ASSIGNMENT_DELAY wci_slvPresent_2$D_IN;
	if (wci_slvPresent_3$EN)
	  wci_slvPresent_3 <= `BSV_ASSIGNMENT_DELAY wci_slvPresent_3$D_IN;
	if (wci_slvPresent_4$EN)
	  wci_slvPresent_4 <= `BSV_ASSIGNMENT_DELAY wci_slvPresent_4$D_IN;
	if (wci_slvPresent_5$EN)
	  wci_slvPresent_5 <= `BSV_ASSIGNMENT_DELAY wci_slvPresent_5$D_IN;
	if (wci_slvPresent_6$EN)
	  wci_slvPresent_6 <= `BSV_ASSIGNMENT_DELAY wci_slvPresent_6$D_IN;
	if (wci_slvPresent_7$EN)
	  wci_slvPresent_7 <= `BSV_ASSIGNMENT_DELAY wci_slvPresent_7$D_IN;
	if (wci_slvPresent_8$EN)
	  wci_slvPresent_8 <= `BSV_ASSIGNMENT_DELAY wci_slvPresent_8$D_IN;
	if (wci_slvPresent_9$EN)
	  wci_slvPresent_9 <= `BSV_ASSIGNMENT_DELAY wci_slvPresent_9$D_IN;
	if (wci_wReset_n$EN)
	  wci_wReset_n <= `BSV_ASSIGNMENT_DELAY wci_wReset_n$D_IN;
	if (wci_wReset_n_1$EN)
	  wci_wReset_n_1 <= `BSV_ASSIGNMENT_DELAY wci_wReset_n_1$D_IN;
	if (wci_wReset_n_10$EN)
	  wci_wReset_n_10 <= `BSV_ASSIGNMENT_DELAY wci_wReset_n_10$D_IN;
	if (wci_wReset_n_11$EN)
	  wci_wReset_n_11 <= `BSV_ASSIGNMENT_DELAY wci_wReset_n_11$D_IN;
	if (wci_wReset_n_12$EN)
	  wci_wReset_n_12 <= `BSV_ASSIGNMENT_DELAY wci_wReset_n_12$D_IN;
	if (wci_wReset_n_13$EN)
	  wci_wReset_n_13 <= `BSV_ASSIGNMENT_DELAY wci_wReset_n_13$D_IN;
	if (wci_wReset_n_14$EN)
	  wci_wReset_n_14 <= `BSV_ASSIGNMENT_DELAY wci_wReset_n_14$D_IN;
	if (wci_wReset_n_2$EN)
	  wci_wReset_n_2 <= `BSV_ASSIGNMENT_DELAY wci_wReset_n_2$D_IN;
	if (wci_wReset_n_3$EN)
	  wci_wReset_n_3 <= `BSV_ASSIGNMENT_DELAY wci_wReset_n_3$D_IN;
	if (wci_wReset_n_4$EN)
	  wci_wReset_n_4 <= `BSV_ASSIGNMENT_DELAY wci_wReset_n_4$D_IN;
	if (wci_wReset_n_5$EN)
	  wci_wReset_n_5 <= `BSV_ASSIGNMENT_DELAY wci_wReset_n_5$D_IN;
	if (wci_wReset_n_6$EN)
	  wci_wReset_n_6 <= `BSV_ASSIGNMENT_DELAY wci_wReset_n_6$D_IN;
	if (wci_wReset_n_7$EN)
	  wci_wReset_n_7 <= `BSV_ASSIGNMENT_DELAY wci_wReset_n_7$D_IN;
	if (wci_wReset_n_8$EN)
	  wci_wReset_n_8 <= `BSV_ASSIGNMENT_DELAY wci_wReset_n_8$D_IN;
	if (wci_wReset_n_9$EN)
	  wci_wReset_n_9 <= `BSV_ASSIGNMENT_DELAY wci_wReset_n_9$D_IN;
	if (wci_wTimeout$EN)
	  wci_wTimeout <= `BSV_ASSIGNMENT_DELAY wci_wTimeout$D_IN;
	if (wci_wTimeout_1$EN)
	  wci_wTimeout_1 <= `BSV_ASSIGNMENT_DELAY wci_wTimeout_1$D_IN;
	if (wci_wTimeout_10$EN)
	  wci_wTimeout_10 <= `BSV_ASSIGNMENT_DELAY wci_wTimeout_10$D_IN;
	if (wci_wTimeout_11$EN)
	  wci_wTimeout_11 <= `BSV_ASSIGNMENT_DELAY wci_wTimeout_11$D_IN;
	if (wci_wTimeout_12$EN)
	  wci_wTimeout_12 <= `BSV_ASSIGNMENT_DELAY wci_wTimeout_12$D_IN;
	if (wci_wTimeout_13$EN)
	  wci_wTimeout_13 <= `BSV_ASSIGNMENT_DELAY wci_wTimeout_13$D_IN;
	if (wci_wTimeout_14$EN)
	  wci_wTimeout_14 <= `BSV_ASSIGNMENT_DELAY wci_wTimeout_14$D_IN;
	if (wci_wTimeout_2$EN)
	  wci_wTimeout_2 <= `BSV_ASSIGNMENT_DELAY wci_wTimeout_2$D_IN;
	if (wci_wTimeout_3$EN)
	  wci_wTimeout_3 <= `BSV_ASSIGNMENT_DELAY wci_wTimeout_3$D_IN;
	if (wci_wTimeout_4$EN)
	  wci_wTimeout_4 <= `BSV_ASSIGNMENT_DELAY wci_wTimeout_4$D_IN;
	if (wci_wTimeout_5$EN)
	  wci_wTimeout_5 <= `BSV_ASSIGNMENT_DELAY wci_wTimeout_5$D_IN;
	if (wci_wTimeout_6$EN)
	  wci_wTimeout_6 <= `BSV_ASSIGNMENT_DELAY wci_wTimeout_6$D_IN;
	if (wci_wTimeout_7$EN)
	  wci_wTimeout_7 <= `BSV_ASSIGNMENT_DELAY wci_wTimeout_7$D_IN;
	if (wci_wTimeout_8$EN)
	  wci_wTimeout_8 <= `BSV_ASSIGNMENT_DELAY wci_wTimeout_8$D_IN;
	if (wci_wTimeout_9$EN)
	  wci_wTimeout_9 <= `BSV_ASSIGNMENT_DELAY wci_wTimeout_9$D_IN;
	if (wrkAct$EN) wrkAct <= `BSV_ASSIGNMENT_DELAY wrkAct$D_IN;
      end
    if (seqTag$EN) seqTag <= `BSV_ASSIGNMENT_DELAY seqTag$D_IN;
`ifdef not
    if (switch_d$EN) switch_d <= `BSV_ASSIGNMENT_DELAY switch_d$D_IN;
`endif
    if (td$EN) td <= `BSV_ASSIGNMENT_DELAY td$D_IN;
    if (wci_wStatus$EN) wci_wStatus <= `BSV_ASSIGNMENT_DELAY wci_wStatus$D_IN;
    if (wci_wStatus_1$EN)
      wci_wStatus_1 <= `BSV_ASSIGNMENT_DELAY wci_wStatus_1$D_IN;
    if (wci_wStatus_10$EN)
      wci_wStatus_10 <= `BSV_ASSIGNMENT_DELAY wci_wStatus_10$D_IN;
    if (wci_wStatus_11$EN)
      wci_wStatus_11 <= `BSV_ASSIGNMENT_DELAY wci_wStatus_11$D_IN;
    if (wci_wStatus_12$EN)
      wci_wStatus_12 <= `BSV_ASSIGNMENT_DELAY wci_wStatus_12$D_IN;
    if (wci_wStatus_13$EN)
      wci_wStatus_13 <= `BSV_ASSIGNMENT_DELAY wci_wStatus_13$D_IN;
    if (wci_wStatus_14$EN)
      wci_wStatus_14 <= `BSV_ASSIGNMENT_DELAY wci_wStatus_14$D_IN;
    if (wci_wStatus_2$EN)
      wci_wStatus_2 <= `BSV_ASSIGNMENT_DELAY wci_wStatus_2$D_IN;
    if (wci_wStatus_3$EN)
      wci_wStatus_3 <= `BSV_ASSIGNMENT_DELAY wci_wStatus_3$D_IN;
    if (wci_wStatus_4$EN)
      wci_wStatus_4 <= `BSV_ASSIGNMENT_DELAY wci_wStatus_4$D_IN;
    if (wci_wStatus_5$EN)
      wci_wStatus_5 <= `BSV_ASSIGNMENT_DELAY wci_wStatus_5$D_IN;
    if (wci_wStatus_6$EN)
      wci_wStatus_6 <= `BSV_ASSIGNMENT_DELAY wci_wStatus_6$D_IN;
    if (wci_wStatus_7$EN)
      wci_wStatus_7 <= `BSV_ASSIGNMENT_DELAY wci_wStatus_7$D_IN;
    if (wci_wStatus_8$EN)
      wci_wStatus_8 <= `BSV_ASSIGNMENT_DELAY wci_wStatus_8$D_IN;
    if (wci_wStatus_9$EN)
      wci_wStatus_9 <= `BSV_ASSIGNMENT_DELAY wci_wStatus_9$D_IN;
  end

`ifdef not
  always@(posedge CLK_time_clk)
  begin
    if (RST_N_time_rst == `BSV_RESET_VALUE)
      begin
        timeServ_delSec <= `BSV_ASSIGNMENT_DELAY 2'd0;
	timeServ_delSecond <= `BSV_ASSIGNMENT_DELAY 50'h1000000000000;
	timeServ_fracInc <= `BSV_ASSIGNMENT_DELAY 50'd1407374;
	timeServ_fracSeconds <= `BSV_ASSIGNMENT_DELAY 50'd0;
	timeServ_jamFrac <= `BSV_ASSIGNMENT_DELAY 1'd0;
	timeServ_jamFracVal <= `BSV_ASSIGNMENT_DELAY 50'd0;
	timeServ_lastSecond <= `BSV_ASSIGNMENT_DELAY 50'd0;
	timeServ_now <= `BSV_ASSIGNMENT_DELAY 64'd0;
	timeServ_ppsDrive <= `BSV_ASSIGNMENT_DELAY 1'd0;
	timeServ_ppsEdgeCount <= `BSV_ASSIGNMENT_DELAY 8'd0;
	timeServ_ppsExtCapture <= `BSV_ASSIGNMENT_DELAY 1'd0;
	timeServ_ppsExtSyncD <= `BSV_ASSIGNMENT_DELAY 1'd0;
	timeServ_ppsExtSync_d1 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	timeServ_ppsExtSync_d2 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	timeServ_ppsLost <= `BSV_ASSIGNMENT_DELAY 1'd0;
	timeServ_ppsOK <= `BSV_ASSIGNMENT_DELAY 1'd0;
	timeServ_refFreeCount <= `BSV_ASSIGNMENT_DELAY 28'd0;
	timeServ_refFreeSamp <= `BSV_ASSIGNMENT_DELAY 28'd0;
	timeServ_refFreeSpan <= `BSV_ASSIGNMENT_DELAY 28'd0;
	timeServ_refFromRise <= `BSV_ASSIGNMENT_DELAY 28'd0;
	timeServ_refPerCount <= `BSV_ASSIGNMENT_DELAY 28'd0;
	timeServ_refSecCount <= `BSV_ASSIGNMENT_DELAY 32'd0;
	timeServ_xo2 <= `BSV_ASSIGNMENT_DELAY 1'd0;
      end
    else
      begin
        if (timeServ_delSec$EN)
	  timeServ_delSec <= `BSV_ASSIGNMENT_DELAY timeServ_delSec$D_IN;
	if (timeServ_delSecond$EN)
	  timeServ_delSecond <= `BSV_ASSIGNMENT_DELAY timeServ_delSecond$D_IN;
	if (timeServ_fracInc$EN)
	  timeServ_fracInc <= `BSV_ASSIGNMENT_DELAY timeServ_fracInc$D_IN;
	if (timeServ_fracSeconds$EN)
	  timeServ_fracSeconds <= `BSV_ASSIGNMENT_DELAY
	      timeServ_fracSeconds$D_IN;
	if (timeServ_jamFrac$EN)
	  timeServ_jamFrac <= `BSV_ASSIGNMENT_DELAY timeServ_jamFrac$D_IN;
	if (timeServ_jamFracVal$EN)
	  timeServ_jamFracVal <= `BSV_ASSIGNMENT_DELAY
	      timeServ_jamFracVal$D_IN;
	if (timeServ_lastSecond$EN)
	  timeServ_lastSecond <= `BSV_ASSIGNMENT_DELAY
	      timeServ_lastSecond$D_IN;
	if (timeServ_now$EN)
	  timeServ_now <= `BSV_ASSIGNMENT_DELAY timeServ_now$D_IN;
	if (timeServ_ppsDrive$EN)
	  timeServ_ppsDrive <= `BSV_ASSIGNMENT_DELAY timeServ_ppsDrive$D_IN;
	if (timeServ_ppsEdgeCount$EN)
	  timeServ_ppsEdgeCount <= `BSV_ASSIGNMENT_DELAY
	      timeServ_ppsEdgeCount$D_IN;
	if (timeServ_ppsExtCapture$EN)
	  timeServ_ppsExtCapture <= `BSV_ASSIGNMENT_DELAY
	      timeServ_ppsExtCapture$D_IN;
	if (timeServ_ppsExtSyncD$EN)
	  timeServ_ppsExtSyncD <= `BSV_ASSIGNMENT_DELAY
	      timeServ_ppsExtSyncD$D_IN;
	if (timeServ_ppsExtSync_d1$EN)
	  timeServ_ppsExtSync_d1 <= `BSV_ASSIGNMENT_DELAY
	      timeServ_ppsExtSync_d1$D_IN;
	if (timeServ_ppsExtSync_d2$EN)
	  timeServ_ppsExtSync_d2 <= `BSV_ASSIGNMENT_DELAY
	      timeServ_ppsExtSync_d2$D_IN;
	if (timeServ_ppsLost$EN)
	  timeServ_ppsLost <= `BSV_ASSIGNMENT_DELAY timeServ_ppsLost$D_IN;
	if (timeServ_ppsOK$EN)
	  timeServ_ppsOK <= `BSV_ASSIGNMENT_DELAY timeServ_ppsOK$D_IN;
	if (timeServ_refFreeCount$EN)
	  timeServ_refFreeCount <= `BSV_ASSIGNMENT_DELAY
	      timeServ_refFreeCount$D_IN;
	if (timeServ_refFreeSamp$EN)
	  timeServ_refFreeSamp <= `BSV_ASSIGNMENT_DELAY
	      timeServ_refFreeSamp$D_IN;
	if (timeServ_refFreeSpan$EN)
	  timeServ_refFreeSpan <= `BSV_ASSIGNMENT_DELAY
	      timeServ_refFreeSpan$D_IN;
	if (timeServ_refFromRise$EN)
	  timeServ_refFromRise <= `BSV_ASSIGNMENT_DELAY
	      timeServ_refFromRise$D_IN;
	if (timeServ_refPerCount$EN)
	  timeServ_refPerCount <= `BSV_ASSIGNMENT_DELAY
	      timeServ_refPerCount$D_IN;
	if (timeServ_refSecCount$EN)
	  timeServ_refSecCount <= `BSV_ASSIGNMENT_DELAY
	      timeServ_refSecCount$D_IN;
	if (timeServ_xo2$EN)
	  timeServ_xo2 <= `BSV_ASSIGNMENT_DELAY timeServ_xo2$D_IN;
      end
  end
`endif

  // synopsys translate_off
  `ifdef BSV_NO_INITIAL_BLOCKS
  `else // not BSV_NO_INITIAL_BLOCKS
  initial
  begin
    cpControl = 32'hAAAAAAAA;
    cpReq = 65'h0AAAAAAAAAAAAAAAA;
`ifdef not
    deltaTime = 64'hAAAAAAAAAAAAAAAA;
`endif
    dispatched = 1'h0;
`ifdef not
    dna_cnt = 7'h2A;
    dna_rdReg = 1'h0;
    dna_shftReg = 1'h0;
    dna_sr = 57'h0AAAAAAAAAAAAAA;
`endif
    readCntReg = 32'hAAAAAAAA;
    rogueTLP = 4'hA;
`ifdef not
    rom_serverAdapter_cnt = 3'h2;
    rom_serverAdapter_s1 = 2'h2;
`endif
    scratch20 = 32'hAAAAAAAA;
    scratch24 = 32'hAAAAAAAA;
    seqTag = 8'hAA;
`ifdef not
    switch_d = 3'h2;
`endif
    td = 32'hAAAAAAAA;
`ifdef not
    timeServ_delSec = 2'h2;
    timeServ_delSecond = 50'h2AAAAAAAAAAAA;
    timeServ_fracInc = 50'h2AAAAAAAAAAAA;
    timeServ_fracSeconds = 50'h2AAAAAAAAAAAA;
    timeServ_gpsInSticky = 1'h0;
    timeServ_jamFrac = 1'h0;
    timeServ_jamFracVal = 50'h2AAAAAAAAAAAA;
    timeServ_lastSecond = 50'h2AAAAAAAAAAAA;
    timeServ_now = 64'hAAAAAAAAAAAAAAAA;
    timeServ_ppsDrive = 1'h0;
    timeServ_ppsEdgeCount = 8'hAA;
    timeServ_ppsExtCapture = 1'h0;
    timeServ_ppsExtSyncD = 1'h0;
    timeServ_ppsExtSync_d1 = 1'h0;
    timeServ_ppsExtSync_d2 = 1'h0;
    timeServ_ppsInSticky = 1'h0;
    timeServ_ppsLost = 1'h0;
    timeServ_ppsLostSticky = 1'h0;
    timeServ_ppsOK = 1'h0;
    timeServ_refFreeCount = 28'hAAAAAAA;
    timeServ_refFreeSamp = 28'hAAAAAAA;
    timeServ_refFreeSpan = 28'hAAAAAAA;
    timeServ_refFromRise = 28'hAAAAAAA;
    timeServ_refPerCount = 28'hAAAAAAA;
    timeServ_refSecCount = 32'hAAAAAAAA;
    timeServ_rplTimeControl = 5'h0A;
    timeServ_timeSetSticky = 1'h0;
    timeServ_xo2 = 1'h0;
`endif
    warmResetP = 1'h0;
    wci_busy = 1'h0;
    wci_busy_1 = 1'h0;
    wci_busy_10 = 1'h0;
    wci_busy_11 = 1'h0;
    wci_busy_12 = 1'h0;
    wci_busy_13 = 1'h0;
    wci_busy_14 = 1'h0;
    wci_busy_2 = 1'h0;
    wci_busy_3 = 1'h0;
    wci_busy_4 = 1'h0;
    wci_busy_5 = 1'h0;
    wci_busy_6 = 1'h0;
    wci_busy_7 = 1'h0;
    wci_busy_8 = 1'h0;
    wci_busy_9 = 1'h0;
    wci_lastConfigAddr = 33'h0AAAAAAAA;
    wci_lastConfigAddr_1 = 33'h0AAAAAAAA;
    wci_lastConfigAddr_10 = 33'h0AAAAAAAA;
    wci_lastConfigAddr_11 = 33'h0AAAAAAAA;
    wci_lastConfigAddr_12 = 33'h0AAAAAAAA;
    wci_lastConfigAddr_13 = 33'h0AAAAAAAA;
    wci_lastConfigAddr_14 = 33'h0AAAAAAAA;
    wci_lastConfigAddr_2 = 33'h0AAAAAAAA;
    wci_lastConfigAddr_3 = 33'h0AAAAAAAA;
    wci_lastConfigAddr_4 = 33'h0AAAAAAAA;
    wci_lastConfigAddr_5 = 33'h0AAAAAAAA;
    wci_lastConfigAddr_6 = 33'h0AAAAAAAA;
    wci_lastConfigAddr_7 = 33'h0AAAAAAAA;
    wci_lastConfigAddr_8 = 33'h0AAAAAAAA;
    wci_lastConfigAddr_9 = 33'h0AAAAAAAA;
    wci_lastConfigBE = 5'h0A;
    wci_lastConfigBE_1 = 5'h0A;
    wci_lastConfigBE_10 = 5'h0A;
    wci_lastConfigBE_11 = 5'h0A;
    wci_lastConfigBE_12 = 5'h0A;
    wci_lastConfigBE_13 = 5'h0A;
    wci_lastConfigBE_14 = 5'h0A;
    wci_lastConfigBE_2 = 5'h0A;
    wci_lastConfigBE_3 = 5'h0A;
    wci_lastConfigBE_4 = 5'h0A;
    wci_lastConfigBE_5 = 5'h0A;
    wci_lastConfigBE_6 = 5'h0A;
    wci_lastConfigBE_7 = 5'h0A;
    wci_lastConfigBE_8 = 5'h0A;
    wci_lastConfigBE_9 = 5'h0A;
    wci_lastControlOp = 4'hA;
    wci_lastControlOp_1 = 4'hA;
    wci_lastControlOp_10 = 4'hA;
    wci_lastControlOp_11 = 4'hA;
    wci_lastControlOp_12 = 4'hA;
    wci_lastControlOp_13 = 4'hA;
    wci_lastControlOp_14 = 4'hA;
    wci_lastControlOp_2 = 4'hA;
    wci_lastControlOp_3 = 4'hA;
    wci_lastControlOp_4 = 4'hA;
    wci_lastControlOp_5 = 4'hA;
    wci_lastControlOp_6 = 4'hA;
    wci_lastControlOp_7 = 4'hA;
    wci_lastControlOp_8 = 4'hA;
    wci_lastControlOp_9 = 4'hA;
    wci_lastOpWrite = 2'h2;
    wci_lastOpWrite_1 = 2'h2;
    wci_lastOpWrite_10 = 2'h2;
    wci_lastOpWrite_11 = 2'h2;
    wci_lastOpWrite_12 = 2'h2;
    wci_lastOpWrite_13 = 2'h2;
    wci_lastOpWrite_14 = 2'h2;
    wci_lastOpWrite_2 = 2'h2;
    wci_lastOpWrite_3 = 2'h2;
    wci_lastOpWrite_4 = 2'h2;
    wci_lastOpWrite_5 = 2'h2;
    wci_lastOpWrite_6 = 2'h2;
    wci_lastOpWrite_7 = 2'h2;
    wci_lastOpWrite_8 = 2'h2;
    wci_lastOpWrite_9 = 2'h2;
    wci_mFlagReg = 2'h2;
    wci_mFlagReg_1 = 2'h2;
    wci_mFlagReg_10 = 2'h2;
    wci_mFlagReg_11 = 2'h2;
    wci_mFlagReg_12 = 2'h2;
    wci_mFlagReg_13 = 2'h2;
    wci_mFlagReg_14 = 2'h2;
    wci_mFlagReg_2 = 2'h2;
    wci_mFlagReg_3 = 2'h2;
    wci_mFlagReg_4 = 2'h2;
    wci_mFlagReg_5 = 2'h2;
    wci_mFlagReg_6 = 2'h2;
    wci_mFlagReg_7 = 2'h2;
    wci_mFlagReg_8 = 2'h2;
    wci_mFlagReg_9 = 2'h2;
    wci_pageWindow = 12'hAAA;
    wci_pageWindow_1 = 12'hAAA;
    wci_pageWindow_10 = 12'hAAA;
    wci_pageWindow_11 = 12'hAAA;
    wci_pageWindow_12 = 12'hAAA;
    wci_pageWindow_13 = 12'hAAA;
    wci_pageWindow_14 = 12'hAAA;
    wci_pageWindow_2 = 12'hAAA;
    wci_pageWindow_3 = 12'hAAA;
    wci_pageWindow_4 = 12'hAAA;
    wci_pageWindow_5 = 12'hAAA;
    wci_pageWindow_6 = 12'hAAA;
    wci_pageWindow_7 = 12'hAAA;
    wci_pageWindow_8 = 12'hAAA;
    wci_pageWindow_9 = 12'hAAA;
    wci_reqERR = 3'h2;
    wci_reqERR_1 = 3'h2;
    wci_reqERR_10 = 3'h2;
    wci_reqERR_11 = 3'h2;
    wci_reqERR_12 = 3'h2;
    wci_reqERR_13 = 3'h2;
    wci_reqERR_14 = 3'h2;
    wci_reqERR_2 = 3'h2;
    wci_reqERR_3 = 3'h2;
    wci_reqERR_4 = 3'h2;
    wci_reqERR_5 = 3'h2;
    wci_reqERR_6 = 3'h2;
    wci_reqERR_7 = 3'h2;
    wci_reqERR_8 = 3'h2;
    wci_reqERR_9 = 3'h2;
    wci_reqFAIL = 3'h2;
    wci_reqFAIL_1 = 3'h2;
    wci_reqFAIL_10 = 3'h2;
    wci_reqFAIL_11 = 3'h2;
    wci_reqFAIL_12 = 3'h2;
    wci_reqFAIL_13 = 3'h2;
    wci_reqFAIL_14 = 3'h2;
    wci_reqFAIL_2 = 3'h2;
    wci_reqFAIL_3 = 3'h2;
    wci_reqFAIL_4 = 3'h2;
    wci_reqFAIL_5 = 3'h2;
    wci_reqFAIL_6 = 3'h2;
    wci_reqFAIL_7 = 3'h2;
    wci_reqFAIL_8 = 3'h2;
    wci_reqFAIL_9 = 3'h2;
    wci_reqF_10_c_r = 1'h0;
    wci_reqF_10_q_0 = 72'hAAAAAAAAAAAAAAAAAA;
    wci_reqF_11_c_r = 1'h0;
    wci_reqF_11_q_0 = 72'hAAAAAAAAAAAAAAAAAA;
    wci_reqF_12_c_r = 1'h0;
    wci_reqF_12_q_0 = 72'hAAAAAAAAAAAAAAAAAA;
    wci_reqF_13_c_r = 1'h0;
    wci_reqF_13_q_0 = 72'hAAAAAAAAAAAAAAAAAA;
    wci_reqF_14_c_r = 1'h0;
    wci_reqF_14_q_0 = 72'hAAAAAAAAAAAAAAAAAA;
    wci_reqF_1_c_r = 1'h0;
    wci_reqF_1_q_0 = 72'hAAAAAAAAAAAAAAAAAA;
    wci_reqF_2_c_r = 1'h0;
    wci_reqF_2_q_0 = 72'hAAAAAAAAAAAAAAAAAA;
    wci_reqF_3_c_r = 1'h0;
    wci_reqF_3_q_0 = 72'hAAAAAAAAAAAAAAAAAA;
    wci_reqF_4_c_r = 1'h0;
    wci_reqF_4_q_0 = 72'hAAAAAAAAAAAAAAAAAA;
    wci_reqF_5_c_r = 1'h0;
    wci_reqF_5_q_0 = 72'hAAAAAAAAAAAAAAAAAA;
    wci_reqF_6_c_r = 1'h0;
    wci_reqF_6_q_0 = 72'hAAAAAAAAAAAAAAAAAA;
    wci_reqF_7_c_r = 1'h0;
    wci_reqF_7_q_0 = 72'hAAAAAAAAAAAAAAAAAA;
    wci_reqF_8_c_r = 1'h0;
    wci_reqF_8_q_0 = 72'hAAAAAAAAAAAAAAAAAA;
    wci_reqF_9_c_r = 1'h0;
    wci_reqF_9_q_0 = 72'hAAAAAAAAAAAAAAAAAA;
    wci_reqF_c_r = 1'h0;
    wci_reqF_q_0 = 72'hAAAAAAAAAAAAAAAAAA;
    wci_reqPend = 2'h2;
    wci_reqPend_1 = 2'h2;
    wci_reqPend_10 = 2'h2;
    wci_reqPend_11 = 2'h2;
    wci_reqPend_12 = 2'h2;
    wci_reqPend_13 = 2'h2;
    wci_reqPend_14 = 2'h2;
    wci_reqPend_2 = 2'h2;
    wci_reqPend_3 = 2'h2;
    wci_reqPend_4 = 2'h2;
    wci_reqPend_5 = 2'h2;
    wci_reqPend_6 = 2'h2;
    wci_reqPend_7 = 2'h2;
    wci_reqPend_8 = 2'h2;
    wci_reqPend_9 = 2'h2;
    wci_reqTO = 3'h2;
    wci_reqTO_1 = 3'h2;
    wci_reqTO_10 = 3'h2;
    wci_reqTO_11 = 3'h2;
    wci_reqTO_12 = 3'h2;
    wci_reqTO_13 = 3'h2;
    wci_reqTO_14 = 3'h2;
    wci_reqTO_2 = 3'h2;
    wci_reqTO_3 = 3'h2;
    wci_reqTO_4 = 3'h2;
    wci_reqTO_5 = 3'h2;
    wci_reqTO_6 = 3'h2;
    wci_reqTO_7 = 3'h2;
    wci_reqTO_8 = 3'h2;
    wci_reqTO_9 = 3'h2;
    wci_respTimr = 32'hAAAAAAAA;
    wci_respTimrAct = 1'h0;
    wci_respTimrAct_1 = 1'h0;
    wci_respTimrAct_10 = 1'h0;
    wci_respTimrAct_11 = 1'h0;
    wci_respTimrAct_12 = 1'h0;
    wci_respTimrAct_13 = 1'h0;
    wci_respTimrAct_14 = 1'h0;
    wci_respTimrAct_2 = 1'h0;
    wci_respTimrAct_3 = 1'h0;
    wci_respTimrAct_4 = 1'h0;
    wci_respTimrAct_5 = 1'h0;
    wci_respTimrAct_6 = 1'h0;
    wci_respTimrAct_7 = 1'h0;
    wci_respTimrAct_8 = 1'h0;
    wci_respTimrAct_9 = 1'h0;
    wci_respTimr_1 = 32'hAAAAAAAA;
    wci_respTimr_10 = 32'hAAAAAAAA;
    wci_respTimr_11 = 32'hAAAAAAAA;
    wci_respTimr_12 = 32'hAAAAAAAA;
    wci_respTimr_13 = 32'hAAAAAAAA;
    wci_respTimr_14 = 32'hAAAAAAAA;
    wci_respTimr_2 = 32'hAAAAAAAA;
    wci_respTimr_3 = 32'hAAAAAAAA;
    wci_respTimr_4 = 32'hAAAAAAAA;
    wci_respTimr_5 = 32'hAAAAAAAA;
    wci_respTimr_6 = 32'hAAAAAAAA;
    wci_respTimr_7 = 32'hAAAAAAAA;
    wci_respTimr_8 = 32'hAAAAAAAA;
    wci_respTimr_9 = 32'hAAAAAAAA;
    wci_sThreadBusy_d = 1'h0;
    wci_sThreadBusy_d_1 = 1'h0;
    wci_sThreadBusy_d_10 = 1'h0;
    wci_sThreadBusy_d_11 = 1'h0;
    wci_sThreadBusy_d_12 = 1'h0;
    wci_sThreadBusy_d_13 = 1'h0;
    wci_sThreadBusy_d_14 = 1'h0;
    wci_sThreadBusy_d_2 = 1'h0;
    wci_sThreadBusy_d_3 = 1'h0;
    wci_sThreadBusy_d_4 = 1'h0;
    wci_sThreadBusy_d_5 = 1'h0;
    wci_sThreadBusy_d_6 = 1'h0;
    wci_sThreadBusy_d_7 = 1'h0;
    wci_sThreadBusy_d_8 = 1'h0;
    wci_sThreadBusy_d_9 = 1'h0;
    wci_sfCap = 1'h0;
    wci_sfCapClear = 1'h0;
    wci_sfCapClear_10 = 1'h0;
    wci_sfCapClear_11 = 1'h0;
    wci_sfCapClear_12 = 1'h0;
    wci_sfCapClear_13 = 1'h0;
    wci_sfCapClear_14 = 1'h0;
    wci_sfCapClear_1_1 = 1'h0;
    wci_sfCapClear_2 = 1'h0;
    wci_sfCapClear_3 = 1'h0;
    wci_sfCapClear_4 = 1'h0;
    wci_sfCapClear_5 = 1'h0;
    wci_sfCapClear_6 = 1'h0;
    wci_sfCapClear_7 = 1'h0;
    wci_sfCapClear_8 = 1'h0;
    wci_sfCapClear_9 = 1'h0;
    wci_sfCapSet = 1'h0;
    wci_sfCapSet_10 = 1'h0;
    wci_sfCapSet_11 = 1'h0;
    wci_sfCapSet_12 = 1'h0;
    wci_sfCapSet_13 = 1'h0;
    wci_sfCapSet_14 = 1'h0;
    wci_sfCapSet_1_1 = 1'h0;
    wci_sfCapSet_2 = 1'h0;
    wci_sfCapSet_3 = 1'h0;
    wci_sfCapSet_4 = 1'h0;
    wci_sfCapSet_5 = 1'h0;
    wci_sfCapSet_6 = 1'h0;
    wci_sfCapSet_7 = 1'h0;
    wci_sfCapSet_8 = 1'h0;
    wci_sfCapSet_9 = 1'h0;
    wci_sfCap_1 = 1'h0;
    wci_sfCap_10 = 1'h0;
    wci_sfCap_11 = 1'h0;
    wci_sfCap_12 = 1'h0;
    wci_sfCap_13 = 1'h0;
    wci_sfCap_14 = 1'h0;
    wci_sfCap_2 = 1'h0;
    wci_sfCap_3 = 1'h0;
    wci_sfCap_4 = 1'h0;
    wci_sfCap_5 = 1'h0;
    wci_sfCap_6 = 1'h0;
    wci_sfCap_7 = 1'h0;
    wci_sfCap_8 = 1'h0;
    wci_sfCap_9 = 1'h0;
    wci_slvPresent = 1'h0;
    wci_slvPresent_1 = 1'h0;
    wci_slvPresent_10 = 1'h0;
    wci_slvPresent_11 = 1'h0;
    wci_slvPresent_12 = 1'h0;
    wci_slvPresent_13 = 1'h0;
    wci_slvPresent_14 = 1'h0;
    wci_slvPresent_2 = 1'h0;
    wci_slvPresent_3 = 1'h0;
    wci_slvPresent_4 = 1'h0;
    wci_slvPresent_5 = 1'h0;
    wci_slvPresent_6 = 1'h0;
    wci_slvPresent_7 = 1'h0;
    wci_slvPresent_8 = 1'h0;
    wci_slvPresent_9 = 1'h0;
    wci_wReset_n = 1'h0;
    wci_wReset_n_1 = 1'h0;
    wci_wReset_n_10 = 1'h0;
    wci_wReset_n_11 = 1'h0;
    wci_wReset_n_12 = 1'h0;
    wci_wReset_n_13 = 1'h0;
    wci_wReset_n_14 = 1'h0;
    wci_wReset_n_2 = 1'h0;
    wci_wReset_n_3 = 1'h0;
    wci_wReset_n_4 = 1'h0;
    wci_wReset_n_5 = 1'h0;
    wci_wReset_n_6 = 1'h0;
    wci_wReset_n_7 = 1'h0;
    wci_wReset_n_8 = 1'h0;
    wci_wReset_n_9 = 1'h0;
    wci_wStatus = 32'hAAAAAAAA;
    wci_wStatus_1 = 32'hAAAAAAAA;
    wci_wStatus_10 = 32'hAAAAAAAA;
    wci_wStatus_11 = 32'hAAAAAAAA;
    wci_wStatus_12 = 32'hAAAAAAAA;
    wci_wStatus_13 = 32'hAAAAAAAA;
    wci_wStatus_14 = 32'hAAAAAAAA;
    wci_wStatus_2 = 32'hAAAAAAAA;
    wci_wStatus_3 = 32'hAAAAAAAA;
    wci_wStatus_4 = 32'hAAAAAAAA;
    wci_wStatus_5 = 32'hAAAAAAAA;
    wci_wStatus_6 = 32'hAAAAAAAA;
    wci_wStatus_7 = 32'hAAAAAAAA;
    wci_wStatus_8 = 32'hAAAAAAAA;
    wci_wStatus_9 = 32'hAAAAAAAA;
    wci_wTimeout = 5'h0A;
    wci_wTimeout_1 = 5'h0A;
    wci_wTimeout_10 = 5'h0A;
    wci_wTimeout_11 = 5'h0A;
    wci_wTimeout_12 = 5'h0A;
    wci_wTimeout_13 = 5'h0A;
    wci_wTimeout_14 = 5'h0A;
    wci_wTimeout_2 = 5'h0A;
    wci_wTimeout_3 = 5'h0A;
    wci_wTimeout_4 = 5'h0A;
    wci_wTimeout_5 = 5'h0A;
    wci_wTimeout_6 = 5'h0A;
    wci_wTimeout_7 = 5'h0A;
    wci_wTimeout_8 = 5'h0A;
    wci_wTimeout_9 = 5'h0A;
    wrkAct = 4'hA;
  end
  `endif // BSV_NO_INITIAL_BLOCKS
  // synopsys translate_on

  // handling of system tasks

  // synopsys translate_off
  always@(negedge CLK)
  begin
    #0;
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_T_T_F)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_T_T_F)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_T_F_T)
	begin
	  v__h79502 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_T_F_T)
	$display("[%0d]: %m: WORKER CONTROL ARM...", v__h79502);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_T_F_T)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_T_F_T)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_T_F_F_F_T)
	begin
	  v__h80094 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_T_F_F_F_T)
	$display("[%0d]: %m: pageWindow register written with %0x ",
		 v__h80094,
		 cpReq[59:28]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_T_F_F_F_T)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_T_F_F_F_T)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_T_F_F_F_F)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_T_F_F_F_F)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_T_T_F)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_T_T_F)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_T_F_T)
	begin
	  v__h80203 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_T_F_T)
	$display("[%0d]: %m: WORKER CONTROL ARM...", v__h80203);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_T_F_T)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_T_F_T)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_T_F_F_F_T)
	begin
	  v__h80782 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_T_F_F_F_T)
	$display("[%0d]: %m: pageWindow register written with %0x ",
		 v__h80782,
		 cpReq[59:28]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_T_F_F_F_T)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_T_F_F_F_T)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_T_F_F_F_F)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_T_F_F_F_F)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_T_F)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_T_F)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_F_T)
	begin
	  v__h80891 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_F_T)
	$display("[%0d]: %m: WORKER CONTROL ARM...", v__h80891);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_F_T)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_F_T)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_F_F_F_T)
	begin
	  v__h81470 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_F_F_F_T)
	$display("[%0d]: %m: pageWindow register written with %0x ",
		 v__h81470,
		 cpReq[59:28]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_F_F_F_T)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_F_F_F_T)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_F_F_F_F)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_F_F_F_F)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_T_F)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_T_F)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_F_T)
	begin
	  v__h81579 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_F_T)
	$display("[%0d]: %m: WORKER CONTROL ARM...", v__h81579);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_F_T)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_F_T)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_F_F_F_T)
	begin
	  v__h82158 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_F_F_F_T)
	$display("[%0d]: %m: pageWindow register written with %0x ",
		 v__h82158,
		 cpReq[59:28]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_F_F_F_T)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_F_F_F_T)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_F_F_F_F)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_F_F_F_F)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_T_F)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_T_F)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_F_T)
	begin
	  v__h82267 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_F_T)
	$display("[%0d]: %m: WORKER CONTROL ARM...", v__h82267);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_F_T)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_F_T)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_F_F_F_T)
	begin
	  v__h82846 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_F_F_F_T)
	$display("[%0d]: %m: pageWindow register written with %0x ",
		 v__h82846,
		 cpReq[59:28]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_F_F_F_T)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_F_F_F_T)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_F_F_F_F)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_F_F_F_F)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_T_F)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_T_F)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_T)
	begin
	  v__h82955 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_T)
	$display("[%0d]: %m: WORKER CONTROL ARM...", v__h82955);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_T)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_T)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_F_F_T)
	begin
	  v__h83534 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_F_F_T)
	$display("[%0d]: %m: pageWindow register written with %0x ",
		 v__h83534,
		 cpReq[59:28]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_F_F_T)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_F_F_T)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_F_F_F)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_F_F_F)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_T_F)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_T_F)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_T)
	begin
	  v__h83643 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_T)
	$display("[%0d]: %m: WORKER CONTROL ARM...", v__h83643);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_T)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_T)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_F_F_T)
	begin
	  v__h84222 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_F_F_T)
	$display("[%0d]: %m: pageWindow register written with %0x ",
		 v__h84222,
		 cpReq[59:28]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_F_F_T)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_F_F_T)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_F_F_F)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_F_F_F)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_T_F)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_T_F)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_T)
	begin
	  v__h84331 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_T)
	$display("[%0d]: %m: WORKER CONTROL ARM...", v__h84331);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_T)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_T)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_F_F_T)
	begin
	  v__h84910 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_F_F_T)
	$display("[%0d]: %m: pageWindow register written with %0x ",
		 v__h84910,
		 cpReq[59:28]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_F_F_T)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_F_F_T)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_F_F_F)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_F_F_F)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_T_F)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_T_F)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_T)
	begin
	  v__h85019 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_T)
	$display("[%0d]: %m: WORKER CONTROL ARM...", v__h85019);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_T)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_T)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_F_F_T)
	begin
	  v__h85598 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_F_F_T)
	$display("[%0d]: %m: pageWindow register written with %0x ",
		 v__h85598,
		 cpReq[59:28]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_F_F_T)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_F_F_T)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_F_F_F)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_F_F_F)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_T_F)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_T_F)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_T)
	begin
	  v__h85707 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_T)
	$display("[%0d]: %m: WORKER CONTROL ARM...", v__h85707);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_T)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_T)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_F_F_T)
	begin
	  v__h86286 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_F_F_T)
	$display("[%0d]: %m: pageWindow register written with %0x ",
		 v__h86286,
		 cpReq[59:28]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_F_F_T)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_F_F_T)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_F_F_F)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_F_F_F)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_T_F)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_T_F)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_T)
	begin
	  v__h86395 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_T)
	$display("[%0d]: %m: WORKER CONTROL ARM...", v__h86395);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_T)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_T)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T)
	begin
	  v__h86974 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T)
	$display("[%0d]: %m: pageWindow register written with %0x ",
		 v__h86974,
		 cpReq[59:28]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_T_F)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_T_F)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_T)
	begin
	  v__h87083 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_T)
	$display("[%0d]: %m: WORKER CONTROL ARM...", v__h87083);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_T)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_T)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T)
	begin
	  v__h87662 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T)
	$display("[%0d]: %m: pageWindow register written with %0x ",
		 v__h87662,
		 cpReq[59:28]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T)
	begin
	  v__h87771 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T)
	$display("[%0d]: %m: WORKER CONTROL ARM...", v__h87771);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T)
	begin
	  v__h88350 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T)
	$display("[%0d]: %m: pageWindow register written with %0x ",
		 v__h88350,
		 cpReq[59:28]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T)
	begin
	  v__h88459 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T)
	$display("[%0d]: %m: WORKER CONTROL ARM...", v__h88459);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T)
	begin
	  v__h89038 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T)
	$display("[%0d]: %m: pageWindow register written with %0x ",
		 v__h89038,
		 cpReq[59:28]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T)
	begin
	  v__h89147 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T)
	$display("[%0d]: %m: WORKER CONTROL ARM...", v__h89147);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T)
	begin
	  v__h89726 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T)
	$display("[%0d]: %m: pageWindow register written with %0x ",
		 v__h89726,
		 cpReq[59:28]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_T_T_F)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_T_T_F)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_T_F_T_F)
	begin
	  v__h97130 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_T_F_T_F)
	$display("[%0d]: %m: WORKER CONTROL ARM...", v__h97130);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_T_F_T_F)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_T_F_T_F)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_T_F_F_T)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_T_F_F_T)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_T_F_F_F_T)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_T_F_F_F_T)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_T_F_F_F_F_T)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_T_F_F_F_F_T)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_T_F_F_F_F_F_T)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_T_F_F_F_F_F_T)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_T_F_F_F_F_F_F)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_T_F_F_F_F_F_F)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_T_F)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_T_F)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_F_T_F)
	begin
	  v__h97202 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_F_T_F)
	$display("[%0d]: %m: WORKER CONTROL ARM...", v__h97202);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_F_T_F)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_F_T_F)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_F_F_T)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_F_F_T)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_F_F_F_T)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_F_F_F_T)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_F_F_F_F_T)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_F_F_F_F_T)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_F_F_F_F_F_T)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_F_F_F_F_F_T)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_F_F_F_F_F_F)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_F_F_F_F_F_F)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_T_F)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_T_F)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_F_T_F)
	begin
	  v__h97274 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_F_T_F)
	$display("[%0d]: %m: WORKER CONTROL ARM...", v__h97274);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_F_T_F)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_F_T_F)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_F_F_T)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_F_F_T)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_F_F_F_T)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_F_F_F_T)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_F_F_F_F_T)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_F_F_F_F_T)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_F_F_F_F_F_T)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_F_F_F_F_F_T)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_F_F_F_F_F_F)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_F_F_F_F_F_F)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_T_F)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_T_F)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_F_T_F)
	begin
	  v__h97346 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_F_T_F)
	$display("[%0d]: %m: WORKER CONTROL ARM...", v__h97346);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_F_T_F)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_F_T_F)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_F_F_T)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_F_F_T)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_F_F_F_T)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_F_F_F_T)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_F_F_F_F_T)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_F_F_F_F_T)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_F_F_F_F_F_T)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_F_F_F_F_F_T)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_F_F_F_F_F_F)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_F_F_F_F_F_F)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_T_F)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_T_F)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_F_T_F)
	begin
	  v__h97418 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_F_T_F)
	$display("[%0d]: %m: WORKER CONTROL ARM...", v__h97418);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_F_T_F)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_F_T_F)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_F_F_T)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_F_F_T)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_F_F_F_T)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_F_F_F_T)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_F_F_F_F_T)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_F_F_F_F_T)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_T_F)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_T_F)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_F_T_F)
	begin
	  v__h97490 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_F_T_F)
	$display("[%0d]: %m: WORKER CONTROL ARM...", v__h97490);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_F_T_F)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_F_T_F)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_F_F_T)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_F_F_T)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_F_F_F_T)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_F_F_F_T)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_T_F)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_T_F)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_F_T_F)
	begin
	  v__h97562 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_F_T_F)
	$display("[%0d]: %m: WORKER CONTROL ARM...", v__h97562);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_F_T_F)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_F_T_F)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_F_F_T)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_F_F_T)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_T_F)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_T_F)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F)
	begin
	  v__h97634 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F)
	$display("[%0d]: %m: WORKER CONTROL ARM...", v__h97634);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F)
	begin
	  v__h97706 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F)
	$display("[%0d]: %m: WORKER CONTROL ARM...", v__h97706);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F)
	begin
	  v__h97778 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F)
	$display("[%0d]: %m: WORKER CONTROL ARM...", v__h97778);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F)
	begin
	  v__h97850 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F)
	$display("[%0d]: %m: WORKER CONTROL ARM...", v__h97850);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F)
	begin
	  v__h97922 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F)
	$display("[%0d]: %m: WORKER CONTROL ARM...", v__h97922);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F)
	begin
	  v__h97994 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F)
	$display("[%0d]: %m: WORKER CONTROL ARM...", v__h97994);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F)
	begin
	  v__h98066 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F)
	$display("[%0d]: %m: WORKER CONTROL ARM...", v__h98066);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_F)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F)
	begin
	  v__h98138 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F)
	$display("[%0d]: %m: WORKER CONTROL ARM...", v__h98138);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_F)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_T)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_T)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_T)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_F_F_F_F)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
`ifdef not
    if (RST_N != `BSV_RESET_VALUE)
      if (rom_serverAdapter_s1[1] && !rom_serverAdapter_outDataCore$FULL_N)
	$display("ERROR: %m: mkBRAMSeverAdapter overrun");
`endif
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_T_F_F_T_T_F)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_T_F_F_T_T_F)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_T_F_F_T_F_F)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_T_F_F_T_F_F)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_T_T_T)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_T_T_T)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_T_F_F_T_T_T)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_T_F_F_T_T_T)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_T_F_F_T_F_T)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_T_F_F_T_F_T)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_T_T_T)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_T_T_T)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_T_F_T_T)
	begin
	  v__h97130 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_T_F_T_T)
	$display("[%0d]: %m: WORKER CONTROL ARM...", v__h97130);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_T_F_T_T)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_T_F_T_T)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_T_F_F_T_T_F)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_T_F_F_T_T_F)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_T_F_F_T_F_F)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_T_F_F_T_F_F)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_T_T_T)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_T_T_T)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_T_F_F_T_T_T)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_T_F_F_T_T_T)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_T_F_F_T_F_T)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_T_F_F_T_F_T)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_T_T)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_T_T)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_F_T_T)
	begin
	  v__h97202 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_F_T_T)
	$display("[%0d]: %m: WORKER CONTROL ARM...", v__h97202);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_F_T_T)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_T_F_T_T)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_F_F_T_T_F)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_F_F_T_T_F)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_F_F_T_F_F)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_F_F_T_F_F)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_T_T)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_T_T)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_F_F_T_T_T)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_F_F_T_T_T)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_F_F_T_F_T)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_T_F_F_T_F_T)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_T_T)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_T_T)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_F_T_T)
	begin
	  v__h97274 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_F_T_T)
	$display("[%0d]: %m: WORKER CONTROL ARM...", v__h97274);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_F_T_T)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_T_F_T_T)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_F_F_T_T_F)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_F_F_T_T_F)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_F_F_T_F_F)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_F_F_T_F_F)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_T_T)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_T_T)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_F_F_T_T_T)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_F_F_T_T_T)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_F_F_T_F_T)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_T_F_F_T_F_T)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_T_T)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_T_T)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_F_T_T)
	begin
	  v__h97346 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_F_T_T)
	$display("[%0d]: %m: WORKER CONTROL ARM...", v__h97346);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_F_T_T)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_T_F_T_T)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_F_F_T_T_F)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_F_F_T_T_F)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_F_F_T_F_F)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_F_F_T_F_F)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_T_T)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_T_T)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_F_F_T_T_T)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_F_F_T_T_T)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_F_F_T_F_T)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_T_F_F_T_F_T)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_T_T)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_T_T)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_F_T_T)
	begin
	  v__h97418 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_F_T_T)
	$display("[%0d]: %m: WORKER CONTROL ARM...", v__h97418);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_F_T_T)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_T_F_T_T)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_F_T_T_F)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_F_T_T_F)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_F_T_F_F)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_F_T_F_F)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_T_T)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_T_T)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_F_T_T_T)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_F_T_T_T)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_F_T_F_T)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_T_F_F_T_F_T)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_T_T)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_T_T)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_F_T_T)
	begin
	  v__h97490 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_F_T_T)
	$display("[%0d]: %m: WORKER CONTROL ARM...", v__h97490);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_F_T_T)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_T_F_T_T)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_F_T_T_F)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_F_T_T_F)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_F_T_F_F)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_F_T_F_F)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_T_T)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_T_T)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_F_T_T_T)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_F_T_T_T)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_F_T_F_T)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_T_F_F_T_F_T)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_T_T)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_T_T)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_F_T_T)
	begin
	  v__h97562 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_F_T_T)
	$display("[%0d]: %m: WORKER CONTROL ARM...", v__h97562);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_F_T_T)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_T_F_T_T)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_F_T_T_F)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_F_T_T_F)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_F_T_F_F)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_F_T_F_F)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_T_T)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_T_T)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_F_T_T_T)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_F_T_T_T)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_F_T_F_T)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_T_F_F_T_F_T)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_T_T)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_T_T)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T)
	begin
	  v__h97634 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T)
	$display("[%0d]: %m: WORKER CONTROL ARM...", v__h97634);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_F_T_T_F)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_F_T_T_F)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_F_T_F_F)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_F_T_F_F)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_T_T)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_T_T)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_F_T_T_T)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_F_T_T_T)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_F_T_F_T)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_T_F_F_T_F_T)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T)
	begin
	  v__h97706 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T)
	$display("[%0d]: %m: WORKER CONTROL ARM...", v__h97706);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_F_T_T_F)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_F_T_T_F)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_F_T_F_F)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_F_T_F_F)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_T_T)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_T_T)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_F_T_F_T)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_T_F_F_T_F_T)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T)
	begin
	  v__h97778 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T)
	$display("[%0d]: %m: WORKER CONTROL ARM...", v__h97778);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_F)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_F)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_F)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_F)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_T_T)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_T_T)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_T)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_T)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T)
	begin
	  v__h97850 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T)
	$display("[%0d]: %m: WORKER CONTROL ARM...", v__h97850);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_F)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_F)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_F)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_F)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_T_T)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_T_T)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_T)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_T)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T)
	begin
	  v__h97922 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T)
	$display("[%0d]: %m: WORKER CONTROL ARM...", v__h97922);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_F)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_F)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_F)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_F)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_T)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_T)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T)
	begin
	  v__h97994 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T)
	$display("[%0d]: %m: WORKER CONTROL ARM...", v__h97994);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_F)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_F)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_F)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_F)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_T)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_T)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T)
	begin
	  v__h98066 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T)
	$display("[%0d]: %m: WORKER CONTROL ARM...", v__h98066);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_F)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_F)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_F)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_F)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_T_T)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_T)
	begin
	  v__h106118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_T_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_F_T_F_T)
	$display("[%0d]: %m: reqWorker WRITE-POSTED   Worker:%0d sp:%x Addr:%0x Data:%0x BE:%0x",
		 v__h106118,
		 _theResult_____1__h76796,
		 cpReq[61:60],
		 cpReq[27:4],
		 cpReq[59:28],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_T_T)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T)
	begin
	  v__h98138 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T)
	$display("[%0d]: %m: WORKER CONTROL ARM...", v__h98138);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T)
	begin
	  v__h106171 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cpDispatch_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_F_T_F_T_T)
	$display("[%0d]: %m: reqWorker READ-REQUESTED Worker:%0d sp:%x Addr:%0x BE:%0x",
		 v__h106171,
		 _theResult_____1__h76814,
		 cpReq[37:36],
		 cpReq[27:4],
		 cpReq[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy && wci_wciResponse$wget[33:32] == 2'd0 &&
	  !wci_respTimr_28_ULT_1_SL_wci_wTimeout_29_30___d5879 &&
	  wci_reqPend == 2'd1)
	begin
	  v__h12057 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy && wci_wciResponse$wget[33:32] == 2'd0 &&
	  !wci_respTimr_28_ULT_1_SL_wci_wTimeout_29_30___d5879 &&
	  wci_reqPend == 2'd1)
	$display("[%0d]: %m: WORKER CONFIG-WRITE TIMEOUT", v__h12057);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy && wci_wciResponse$wget[33:32] == 2'd0 &&
	  !wci_respTimr_28_ULT_1_SL_wci_wTimeout_29_30___d5879 &&
	  wci_reqPend == 2'd2)
	begin
	  v__h12147 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy && wci_wciResponse$wget[33:32] == 2'd0 &&
	  !wci_respTimr_28_ULT_1_SL_wci_wTimeout_29_30___d5879 &&
	  wci_reqPend == 2'd2)
	$display("[%0d]: %m: WORKER CONFIG-READ  TIMEOUT", v__h12147);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy && wci_wciResponse$wget[33:32] == 2'd0 &&
	  !wci_respTimr_28_ULT_1_SL_wci_wTimeout_29_30___d5879 &&
	  wci_reqPend == 2'd3)
	begin
	  v__h12236 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy && wci_wciResponse$wget[33:32] == 2'd0 &&
	  !wci_respTimr_28_ULT_1_SL_wci_wTimeout_29_30___d5879 &&
	  wci_reqPend == 2'd3)
	$display("[%0d]: %m: WORKER CONTROL-OP   TIMEOUT", v__h12236);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy && wci_wciResponse$wget[33:32] == 2'd2 &&
	  wci_reqPend == 2'd1)
	begin
	  v__h12460 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy && wci_wciResponse$wget[33:32] == 2'd2 &&
	  wci_reqPend == 2'd1)
	$display("[%0d]: %m: WORKER CONFIG-WRITE RESPONSE-FAIL", v__h12460);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy && wci_wciResponse$wget[33:32] == 2'd2 &&
	  wci_reqPend == 2'd2)
	begin
	  v__h12550 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy && wci_wciResponse$wget[33:32] == 2'd2 &&
	  wci_reqPend == 2'd2)
	$display("[%0d]: %m: WORKER CONFIG-READ  RESPONSE-FAIL", v__h12550);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy && wci_wciResponse$wget[33:32] == 2'd2 &&
	  wci_reqPend == 2'd3)
	begin
	  v__h12639 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy && wci_wciResponse$wget[33:32] == 2'd2 &&
	  wci_reqPend == 2'd3)
	$display("[%0d]: %m: WORKER CONTROL-OP   RESPONSE-FAIL", v__h12639);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy && wci_wciResponse$wget[33:32] == 2'd3 &&
	  wci_reqPend == 2'd1)
	begin
	  v__h12868 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy && wci_wciResponse$wget[33:32] == 2'd3 &&
	  wci_reqPend == 2'd1)
	$display("[%0d]: %m: WORKER CONFIG-WRITE RESPONSE-ERR", v__h12868);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy && wci_wciResponse$wget[33:32] == 2'd3 &&
	  wci_reqPend == 2'd2)
	begin
	  v__h12958 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy && wci_wciResponse$wget[33:32] == 2'd3 &&
	  wci_reqPend == 2'd2)
	$display("[%0d]: %m: WORKER CONFIG-READ  RESPONSE-ERR", v__h12958);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy && wci_wciResponse$wget[33:32] == 2'd3 &&
	  wci_reqPend == 2'd3)
	begin
	  v__h13047 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy && wci_wciResponse$wget[33:32] == 2'd3 &&
	  wci_reqPend == 2'd3)
	$display("[%0d]: %m: WORKER CONTROL-OP   RESPONSE-ERR", v__h13047);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_1 &&
	  wci_wciResponse_1$wget[33:32] == 2'd0 &&
	  !wci_respTimr_1_68_ULT_1_SL_wci_wTimeout_1_69_70___d5880 &&
	  wci_reqPend_1 == 2'd1)
	begin
	  v__h16497 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_1 &&
	  wci_wciResponse_1$wget[33:32] == 2'd0 &&
	  !wci_respTimr_1_68_ULT_1_SL_wci_wTimeout_1_69_70___d5880 &&
	  wci_reqPend_1 == 2'd1)
	$display("[%0d]: %m: WORKER CONFIG-WRITE TIMEOUT", v__h16497);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_1 &&
	  wci_wciResponse_1$wget[33:32] == 2'd0 &&
	  !wci_respTimr_1_68_ULT_1_SL_wci_wTimeout_1_69_70___d5880 &&
	  wci_reqPend_1 == 2'd2)
	begin
	  v__h16587 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_1 &&
	  wci_wciResponse_1$wget[33:32] == 2'd0 &&
	  !wci_respTimr_1_68_ULT_1_SL_wci_wTimeout_1_69_70___d5880 &&
	  wci_reqPend_1 == 2'd2)
	$display("[%0d]: %m: WORKER CONFIG-READ  TIMEOUT", v__h16587);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_1 &&
	  wci_wciResponse_1$wget[33:32] == 2'd0 &&
	  !wci_respTimr_1_68_ULT_1_SL_wci_wTimeout_1_69_70___d5880 &&
	  wci_reqPend_1 == 2'd3)
	begin
	  v__h16676 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_1 &&
	  wci_wciResponse_1$wget[33:32] == 2'd0 &&
	  !wci_respTimr_1_68_ULT_1_SL_wci_wTimeout_1_69_70___d5880 &&
	  wci_reqPend_1 == 2'd3)
	$display("[%0d]: %m: WORKER CONTROL-OP   TIMEOUT", v__h16676);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_1 &&
	  wci_wciResponse_1$wget[33:32] == 2'd2 &&
	  wci_reqPend_1 == 2'd1)
	begin
	  v__h16900 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_1 &&
	  wci_wciResponse_1$wget[33:32] == 2'd2 &&
	  wci_reqPend_1 == 2'd1)
	$display("[%0d]: %m: WORKER CONFIG-WRITE RESPONSE-FAIL", v__h16900);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_1 &&
	  wci_wciResponse_1$wget[33:32] == 2'd2 &&
	  wci_reqPend_1 == 2'd2)
	begin
	  v__h16990 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_1 &&
	  wci_wciResponse_1$wget[33:32] == 2'd2 &&
	  wci_reqPend_1 == 2'd2)
	$display("[%0d]: %m: WORKER CONFIG-READ  RESPONSE-FAIL", v__h16990);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_1 &&
	  wci_wciResponse_1$wget[33:32] == 2'd2 &&
	  wci_reqPend_1 == 2'd3)
	begin
	  v__h17079 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_1 &&
	  wci_wciResponse_1$wget[33:32] == 2'd2 &&
	  wci_reqPend_1 == 2'd3)
	$display("[%0d]: %m: WORKER CONTROL-OP   RESPONSE-FAIL", v__h17079);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_1 &&
	  wci_wciResponse_1$wget[33:32] == 2'd3 &&
	  wci_reqPend_1 == 2'd1)
	begin
	  v__h17308 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_1 &&
	  wci_wciResponse_1$wget[33:32] == 2'd3 &&
	  wci_reqPend_1 == 2'd1)
	$display("[%0d]: %m: WORKER CONFIG-WRITE RESPONSE-ERR", v__h17308);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_1 &&
	  wci_wciResponse_1$wget[33:32] == 2'd3 &&
	  wci_reqPend_1 == 2'd2)
	begin
	  v__h17398 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_1 &&
	  wci_wciResponse_1$wget[33:32] == 2'd3 &&
	  wci_reqPend_1 == 2'd2)
	$display("[%0d]: %m: WORKER CONFIG-READ  RESPONSE-ERR", v__h17398);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_1 &&
	  wci_wciResponse_1$wget[33:32] == 2'd3 &&
	  wci_reqPend_1 == 2'd3)
	begin
	  v__h17487 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_1 &&
	  wci_wciResponse_1$wget[33:32] == 2'd3 &&
	  wci_reqPend_1 == 2'd3)
	$display("[%0d]: %m: WORKER CONTROL-OP   RESPONSE-ERR", v__h17487);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_2 &&
	  wci_wciResponse_2$wget[33:32] == 2'd0 &&
	  !wci_respTimr_2_08_ULT_1_SL_wci_wTimeout_2_09_10___d5881 &&
	  wci_reqPend_2 == 2'd1)
	begin
	  v__h20937 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_2 &&
	  wci_wciResponse_2$wget[33:32] == 2'd0 &&
	  !wci_respTimr_2_08_ULT_1_SL_wci_wTimeout_2_09_10___d5881 &&
	  wci_reqPend_2 == 2'd1)
	$display("[%0d]: %m: WORKER CONFIG-WRITE TIMEOUT", v__h20937);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_2 &&
	  wci_wciResponse_2$wget[33:32] == 2'd0 &&
	  !wci_respTimr_2_08_ULT_1_SL_wci_wTimeout_2_09_10___d5881 &&
	  wci_reqPend_2 == 2'd2)
	begin
	  v__h21027 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_2 &&
	  wci_wciResponse_2$wget[33:32] == 2'd0 &&
	  !wci_respTimr_2_08_ULT_1_SL_wci_wTimeout_2_09_10___d5881 &&
	  wci_reqPend_2 == 2'd2)
	$display("[%0d]: %m: WORKER CONFIG-READ  TIMEOUT", v__h21027);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_2 &&
	  wci_wciResponse_2$wget[33:32] == 2'd0 &&
	  !wci_respTimr_2_08_ULT_1_SL_wci_wTimeout_2_09_10___d5881 &&
	  wci_reqPend_2 == 2'd3)
	begin
	  v__h21116 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_2 &&
	  wci_wciResponse_2$wget[33:32] == 2'd0 &&
	  !wci_respTimr_2_08_ULT_1_SL_wci_wTimeout_2_09_10___d5881 &&
	  wci_reqPend_2 == 2'd3)
	$display("[%0d]: %m: WORKER CONTROL-OP   TIMEOUT", v__h21116);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_2 &&
	  wci_wciResponse_2$wget[33:32] == 2'd2 &&
	  wci_reqPend_2 == 2'd1)
	begin
	  v__h21340 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_2 &&
	  wci_wciResponse_2$wget[33:32] == 2'd2 &&
	  wci_reqPend_2 == 2'd1)
	$display("[%0d]: %m: WORKER CONFIG-WRITE RESPONSE-FAIL", v__h21340);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_2 &&
	  wci_wciResponse_2$wget[33:32] == 2'd2 &&
	  wci_reqPend_2 == 2'd2)
	begin
	  v__h21430 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_2 &&
	  wci_wciResponse_2$wget[33:32] == 2'd2 &&
	  wci_reqPend_2 == 2'd2)
	$display("[%0d]: %m: WORKER CONFIG-READ  RESPONSE-FAIL", v__h21430);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_2 &&
	  wci_wciResponse_2$wget[33:32] == 2'd2 &&
	  wci_reqPend_2 == 2'd3)
	begin
	  v__h21519 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_2 &&
	  wci_wciResponse_2$wget[33:32] == 2'd2 &&
	  wci_reqPend_2 == 2'd3)
	$display("[%0d]: %m: WORKER CONTROL-OP   RESPONSE-FAIL", v__h21519);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_2 &&
	  wci_wciResponse_2$wget[33:32] == 2'd3 &&
	  wci_reqPend_2 == 2'd1)
	begin
	  v__h21748 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_2 &&
	  wci_wciResponse_2$wget[33:32] == 2'd3 &&
	  wci_reqPend_2 == 2'd1)
	$display("[%0d]: %m: WORKER CONFIG-WRITE RESPONSE-ERR", v__h21748);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_2 &&
	  wci_wciResponse_2$wget[33:32] == 2'd3 &&
	  wci_reqPend_2 == 2'd2)
	begin
	  v__h21838 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_2 &&
	  wci_wciResponse_2$wget[33:32] == 2'd3 &&
	  wci_reqPend_2 == 2'd2)
	$display("[%0d]: %m: WORKER CONFIG-READ  RESPONSE-ERR", v__h21838);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_2 &&
	  wci_wciResponse_2$wget[33:32] == 2'd3 &&
	  wci_reqPend_2 == 2'd3)
	begin
	  v__h21927 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_2 &&
	  wci_wciResponse_2$wget[33:32] == 2'd3 &&
	  wci_reqPend_2 == 2'd3)
	$display("[%0d]: %m: WORKER CONTROL-OP   RESPONSE-ERR", v__h21927);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_3 &&
	  wci_wciResponse_3$wget[33:32] == 2'd0 &&
	  !wci_respTimr_3_48_ULT_1_SL_wci_wTimeout_3_49_50___d5882 &&
	  wci_reqPend_3 == 2'd1)
	begin
	  v__h25377 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_3 &&
	  wci_wciResponse_3$wget[33:32] == 2'd0 &&
	  !wci_respTimr_3_48_ULT_1_SL_wci_wTimeout_3_49_50___d5882 &&
	  wci_reqPend_3 == 2'd1)
	$display("[%0d]: %m: WORKER CONFIG-WRITE TIMEOUT", v__h25377);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_3 &&
	  wci_wciResponse_3$wget[33:32] == 2'd0 &&
	  !wci_respTimr_3_48_ULT_1_SL_wci_wTimeout_3_49_50___d5882 &&
	  wci_reqPend_3 == 2'd2)
	begin
	  v__h25467 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_3 &&
	  wci_wciResponse_3$wget[33:32] == 2'd0 &&
	  !wci_respTimr_3_48_ULT_1_SL_wci_wTimeout_3_49_50___d5882 &&
	  wci_reqPend_3 == 2'd2)
	$display("[%0d]: %m: WORKER CONFIG-READ  TIMEOUT", v__h25467);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_3 &&
	  wci_wciResponse_3$wget[33:32] == 2'd0 &&
	  !wci_respTimr_3_48_ULT_1_SL_wci_wTimeout_3_49_50___d5882 &&
	  wci_reqPend_3 == 2'd3)
	begin
	  v__h25556 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_3 &&
	  wci_wciResponse_3$wget[33:32] == 2'd0 &&
	  !wci_respTimr_3_48_ULT_1_SL_wci_wTimeout_3_49_50___d5882 &&
	  wci_reqPend_3 == 2'd3)
	$display("[%0d]: %m: WORKER CONTROL-OP   TIMEOUT", v__h25556);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_3 &&
	  wci_wciResponse_3$wget[33:32] == 2'd2 &&
	  wci_reqPend_3 == 2'd1)
	begin
	  v__h25780 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_3 &&
	  wci_wciResponse_3$wget[33:32] == 2'd2 &&
	  wci_reqPend_3 == 2'd1)
	$display("[%0d]: %m: WORKER CONFIG-WRITE RESPONSE-FAIL", v__h25780);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_3 &&
	  wci_wciResponse_3$wget[33:32] == 2'd2 &&
	  wci_reqPend_3 == 2'd2)
	begin
	  v__h25870 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_3 &&
	  wci_wciResponse_3$wget[33:32] == 2'd2 &&
	  wci_reqPend_3 == 2'd2)
	$display("[%0d]: %m: WORKER CONFIG-READ  RESPONSE-FAIL", v__h25870);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_3 &&
	  wci_wciResponse_3$wget[33:32] == 2'd2 &&
	  wci_reqPend_3 == 2'd3)
	begin
	  v__h25959 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_3 &&
	  wci_wciResponse_3$wget[33:32] == 2'd2 &&
	  wci_reqPend_3 == 2'd3)
	$display("[%0d]: %m: WORKER CONTROL-OP   RESPONSE-FAIL", v__h25959);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_3 &&
	  wci_wciResponse_3$wget[33:32] == 2'd3 &&
	  wci_reqPend_3 == 2'd1)
	begin
	  v__h26188 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_3 &&
	  wci_wciResponse_3$wget[33:32] == 2'd3 &&
	  wci_reqPend_3 == 2'd1)
	$display("[%0d]: %m: WORKER CONFIG-WRITE RESPONSE-ERR", v__h26188);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_3 &&
	  wci_wciResponse_3$wget[33:32] == 2'd3 &&
	  wci_reqPend_3 == 2'd2)
	begin
	  v__h26278 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_3 &&
	  wci_wciResponse_3$wget[33:32] == 2'd3 &&
	  wci_reqPend_3 == 2'd2)
	$display("[%0d]: %m: WORKER CONFIG-READ  RESPONSE-ERR", v__h26278);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_3 &&
	  wci_wciResponse_3$wget[33:32] == 2'd3 &&
	  wci_reqPend_3 == 2'd3)
	begin
	  v__h26367 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_3 &&
	  wci_wciResponse_3$wget[33:32] == 2'd3 &&
	  wci_reqPend_3 == 2'd3)
	$display("[%0d]: %m: WORKER CONTROL-OP   RESPONSE-ERR", v__h26367);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_4 &&
	  wci_wciResponse_4$wget[33:32] == 2'd0 &&
	  !wci_respTimr_4_88_ULT_1_SL_wci_wTimeout_4_89_90___d5883 &&
	  wci_reqPend_4 == 2'd1)
	begin
	  v__h29817 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_4 &&
	  wci_wciResponse_4$wget[33:32] == 2'd0 &&
	  !wci_respTimr_4_88_ULT_1_SL_wci_wTimeout_4_89_90___d5883 &&
	  wci_reqPend_4 == 2'd1)
	$display("[%0d]: %m: WORKER CONFIG-WRITE TIMEOUT", v__h29817);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_4 &&
	  wci_wciResponse_4$wget[33:32] == 2'd0 &&
	  !wci_respTimr_4_88_ULT_1_SL_wci_wTimeout_4_89_90___d5883 &&
	  wci_reqPend_4 == 2'd2)
	begin
	  v__h29907 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_4 &&
	  wci_wciResponse_4$wget[33:32] == 2'd0 &&
	  !wci_respTimr_4_88_ULT_1_SL_wci_wTimeout_4_89_90___d5883 &&
	  wci_reqPend_4 == 2'd2)
	$display("[%0d]: %m: WORKER CONFIG-READ  TIMEOUT", v__h29907);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_4 &&
	  wci_wciResponse_4$wget[33:32] == 2'd0 &&
	  !wci_respTimr_4_88_ULT_1_SL_wci_wTimeout_4_89_90___d5883 &&
	  wci_reqPend_4 == 2'd3)
	begin
	  v__h29996 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_4 &&
	  wci_wciResponse_4$wget[33:32] == 2'd0 &&
	  !wci_respTimr_4_88_ULT_1_SL_wci_wTimeout_4_89_90___d5883 &&
	  wci_reqPend_4 == 2'd3)
	$display("[%0d]: %m: WORKER CONTROL-OP   TIMEOUT", v__h29996);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_4 &&
	  wci_wciResponse_4$wget[33:32] == 2'd2 &&
	  wci_reqPend_4 == 2'd1)
	begin
	  v__h30220 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_4 &&
	  wci_wciResponse_4$wget[33:32] == 2'd2 &&
	  wci_reqPend_4 == 2'd1)
	$display("[%0d]: %m: WORKER CONFIG-WRITE RESPONSE-FAIL", v__h30220);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_4 &&
	  wci_wciResponse_4$wget[33:32] == 2'd2 &&
	  wci_reqPend_4 == 2'd2)
	begin
	  v__h30310 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_4 &&
	  wci_wciResponse_4$wget[33:32] == 2'd2 &&
	  wci_reqPend_4 == 2'd2)
	$display("[%0d]: %m: WORKER CONFIG-READ  RESPONSE-FAIL", v__h30310);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_4 &&
	  wci_wciResponse_4$wget[33:32] == 2'd2 &&
	  wci_reqPend_4 == 2'd3)
	begin
	  v__h30399 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_4 &&
	  wci_wciResponse_4$wget[33:32] == 2'd2 &&
	  wci_reqPend_4 == 2'd3)
	$display("[%0d]: %m: WORKER CONTROL-OP   RESPONSE-FAIL", v__h30399);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_4 &&
	  wci_wciResponse_4$wget[33:32] == 2'd3 &&
	  wci_reqPend_4 == 2'd1)
	begin
	  v__h30628 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_4 &&
	  wci_wciResponse_4$wget[33:32] == 2'd3 &&
	  wci_reqPend_4 == 2'd1)
	$display("[%0d]: %m: WORKER CONFIG-WRITE RESPONSE-ERR", v__h30628);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_4 &&
	  wci_wciResponse_4$wget[33:32] == 2'd3 &&
	  wci_reqPend_4 == 2'd2)
	begin
	  v__h30718 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_4 &&
	  wci_wciResponse_4$wget[33:32] == 2'd3 &&
	  wci_reqPend_4 == 2'd2)
	$display("[%0d]: %m: WORKER CONFIG-READ  RESPONSE-ERR", v__h30718);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_4 &&
	  wci_wciResponse_4$wget[33:32] == 2'd3 &&
	  wci_reqPend_4 == 2'd3)
	begin
	  v__h30807 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_4 &&
	  wci_wciResponse_4$wget[33:32] == 2'd3 &&
	  wci_reqPend_4 == 2'd3)
	$display("[%0d]: %m: WORKER CONTROL-OP   RESPONSE-ERR", v__h30807);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_5 &&
	  wci_wciResponse_5$wget[33:32] == 2'd0 &&
	  !wci_respTimr_5_28_ULT_1_SL_wci_wTimeout_5_29_30___d5884 &&
	  wci_reqPend_5 == 2'd1)
	begin
	  v__h34257 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_5 &&
	  wci_wciResponse_5$wget[33:32] == 2'd0 &&
	  !wci_respTimr_5_28_ULT_1_SL_wci_wTimeout_5_29_30___d5884 &&
	  wci_reqPend_5 == 2'd1)
	$display("[%0d]: %m: WORKER CONFIG-WRITE TIMEOUT", v__h34257);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_5 &&
	  wci_wciResponse_5$wget[33:32] == 2'd0 &&
	  !wci_respTimr_5_28_ULT_1_SL_wci_wTimeout_5_29_30___d5884 &&
	  wci_reqPend_5 == 2'd2)
	begin
	  v__h34347 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_5 &&
	  wci_wciResponse_5$wget[33:32] == 2'd0 &&
	  !wci_respTimr_5_28_ULT_1_SL_wci_wTimeout_5_29_30___d5884 &&
	  wci_reqPend_5 == 2'd2)
	$display("[%0d]: %m: WORKER CONFIG-READ  TIMEOUT", v__h34347);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_5 &&
	  wci_wciResponse_5$wget[33:32] == 2'd0 &&
	  !wci_respTimr_5_28_ULT_1_SL_wci_wTimeout_5_29_30___d5884 &&
	  wci_reqPend_5 == 2'd3)
	begin
	  v__h34436 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_5 &&
	  wci_wciResponse_5$wget[33:32] == 2'd0 &&
	  !wci_respTimr_5_28_ULT_1_SL_wci_wTimeout_5_29_30___d5884 &&
	  wci_reqPend_5 == 2'd3)
	$display("[%0d]: %m: WORKER CONTROL-OP   TIMEOUT", v__h34436);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_5 &&
	  wci_wciResponse_5$wget[33:32] == 2'd2 &&
	  wci_reqPend_5 == 2'd1)
	begin
	  v__h34660 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_5 &&
	  wci_wciResponse_5$wget[33:32] == 2'd2 &&
	  wci_reqPend_5 == 2'd1)
	$display("[%0d]: %m: WORKER CONFIG-WRITE RESPONSE-FAIL", v__h34660);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_5 &&
	  wci_wciResponse_5$wget[33:32] == 2'd2 &&
	  wci_reqPend_5 == 2'd2)
	begin
	  v__h34750 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_5 &&
	  wci_wciResponse_5$wget[33:32] == 2'd2 &&
	  wci_reqPend_5 == 2'd2)
	$display("[%0d]: %m: WORKER CONFIG-READ  RESPONSE-FAIL", v__h34750);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_5 &&
	  wci_wciResponse_5$wget[33:32] == 2'd2 &&
	  wci_reqPend_5 == 2'd3)
	begin
	  v__h34839 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_5 &&
	  wci_wciResponse_5$wget[33:32] == 2'd2 &&
	  wci_reqPend_5 == 2'd3)
	$display("[%0d]: %m: WORKER CONTROL-OP   RESPONSE-FAIL", v__h34839);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_5 &&
	  wci_wciResponse_5$wget[33:32] == 2'd3 &&
	  wci_reqPend_5 == 2'd1)
	begin
	  v__h35068 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_5 &&
	  wci_wciResponse_5$wget[33:32] == 2'd3 &&
	  wci_reqPend_5 == 2'd1)
	$display("[%0d]: %m: WORKER CONFIG-WRITE RESPONSE-ERR", v__h35068);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_5 &&
	  wci_wciResponse_5$wget[33:32] == 2'd3 &&
	  wci_reqPend_5 == 2'd2)
	begin
	  v__h35158 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_5 &&
	  wci_wciResponse_5$wget[33:32] == 2'd3 &&
	  wci_reqPend_5 == 2'd2)
	$display("[%0d]: %m: WORKER CONFIG-READ  RESPONSE-ERR", v__h35158);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_5 &&
	  wci_wciResponse_5$wget[33:32] == 2'd3 &&
	  wci_reqPend_5 == 2'd3)
	begin
	  v__h35247 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_5 &&
	  wci_wciResponse_5$wget[33:32] == 2'd3 &&
	  wci_reqPend_5 == 2'd3)
	$display("[%0d]: %m: WORKER CONTROL-OP   RESPONSE-ERR", v__h35247);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_6 &&
	  wci_wciResponse_6$wget[33:32] == 2'd0 &&
	  !wci_respTimr_6_068_ULT_1_SL_wci_wTimeout_6_069_ETC___d5885 &&
	  wci_reqPend_6 == 2'd1)
	begin
	  v__h38697 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_6 &&
	  wci_wciResponse_6$wget[33:32] == 2'd0 &&
	  !wci_respTimr_6_068_ULT_1_SL_wci_wTimeout_6_069_ETC___d5885 &&
	  wci_reqPend_6 == 2'd1)
	$display("[%0d]: %m: WORKER CONFIG-WRITE TIMEOUT", v__h38697);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_6 &&
	  wci_wciResponse_6$wget[33:32] == 2'd0 &&
	  !wci_respTimr_6_068_ULT_1_SL_wci_wTimeout_6_069_ETC___d5885 &&
	  wci_reqPend_6 == 2'd2)
	begin
	  v__h38787 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_6 &&
	  wci_wciResponse_6$wget[33:32] == 2'd0 &&
	  !wci_respTimr_6_068_ULT_1_SL_wci_wTimeout_6_069_ETC___d5885 &&
	  wci_reqPend_6 == 2'd2)
	$display("[%0d]: %m: WORKER CONFIG-READ  TIMEOUT", v__h38787);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_6 &&
	  wci_wciResponse_6$wget[33:32] == 2'd0 &&
	  !wci_respTimr_6_068_ULT_1_SL_wci_wTimeout_6_069_ETC___d5885 &&
	  wci_reqPend_6 == 2'd3)
	begin
	  v__h38876 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_6 &&
	  wci_wciResponse_6$wget[33:32] == 2'd0 &&
	  !wci_respTimr_6_068_ULT_1_SL_wci_wTimeout_6_069_ETC___d5885 &&
	  wci_reqPend_6 == 2'd3)
	$display("[%0d]: %m: WORKER CONTROL-OP   TIMEOUT", v__h38876);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_6 &&
	  wci_wciResponse_6$wget[33:32] == 2'd2 &&
	  wci_reqPend_6 == 2'd1)
	begin
	  v__h39100 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_6 &&
	  wci_wciResponse_6$wget[33:32] == 2'd2 &&
	  wci_reqPend_6 == 2'd1)
	$display("[%0d]: %m: WORKER CONFIG-WRITE RESPONSE-FAIL", v__h39100);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_6 &&
	  wci_wciResponse_6$wget[33:32] == 2'd2 &&
	  wci_reqPend_6 == 2'd2)
	begin
	  v__h39190 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_6 &&
	  wci_wciResponse_6$wget[33:32] == 2'd2 &&
	  wci_reqPend_6 == 2'd2)
	$display("[%0d]: %m: WORKER CONFIG-READ  RESPONSE-FAIL", v__h39190);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_6 &&
	  wci_wciResponse_6$wget[33:32] == 2'd2 &&
	  wci_reqPend_6 == 2'd3)
	begin
	  v__h39279 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_6 &&
	  wci_wciResponse_6$wget[33:32] == 2'd2 &&
	  wci_reqPend_6 == 2'd3)
	$display("[%0d]: %m: WORKER CONTROL-OP   RESPONSE-FAIL", v__h39279);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_6 &&
	  wci_wciResponse_6$wget[33:32] == 2'd3 &&
	  wci_reqPend_6 == 2'd1)
	begin
	  v__h39508 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_6 &&
	  wci_wciResponse_6$wget[33:32] == 2'd3 &&
	  wci_reqPend_6 == 2'd1)
	$display("[%0d]: %m: WORKER CONFIG-WRITE RESPONSE-ERR", v__h39508);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_6 &&
	  wci_wciResponse_6$wget[33:32] == 2'd3 &&
	  wci_reqPend_6 == 2'd2)
	begin
	  v__h39598 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_6 &&
	  wci_wciResponse_6$wget[33:32] == 2'd3 &&
	  wci_reqPend_6 == 2'd2)
	$display("[%0d]: %m: WORKER CONFIG-READ  RESPONSE-ERR", v__h39598);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_6 &&
	  wci_wciResponse_6$wget[33:32] == 2'd3 &&
	  wci_reqPend_6 == 2'd3)
	begin
	  v__h39687 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_6 &&
	  wci_wciResponse_6$wget[33:32] == 2'd3 &&
	  wci_reqPend_6 == 2'd3)
	$display("[%0d]: %m: WORKER CONTROL-OP   RESPONSE-ERR", v__h39687);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_7 &&
	  wci_wciResponse_7$wget[33:32] == 2'd0 &&
	  !wci_respTimr_7_208_ULT_1_SL_wci_wTimeout_7_209_ETC___d5886 &&
	  wci_reqPend_7 == 2'd1)
	begin
	  v__h43137 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_7 &&
	  wci_wciResponse_7$wget[33:32] == 2'd0 &&
	  !wci_respTimr_7_208_ULT_1_SL_wci_wTimeout_7_209_ETC___d5886 &&
	  wci_reqPend_7 == 2'd1)
	$display("[%0d]: %m: WORKER CONFIG-WRITE TIMEOUT", v__h43137);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_7 &&
	  wci_wciResponse_7$wget[33:32] == 2'd0 &&
	  !wci_respTimr_7_208_ULT_1_SL_wci_wTimeout_7_209_ETC___d5886 &&
	  wci_reqPend_7 == 2'd2)
	begin
	  v__h43227 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_7 &&
	  wci_wciResponse_7$wget[33:32] == 2'd0 &&
	  !wci_respTimr_7_208_ULT_1_SL_wci_wTimeout_7_209_ETC___d5886 &&
	  wci_reqPend_7 == 2'd2)
	$display("[%0d]: %m: WORKER CONFIG-READ  TIMEOUT", v__h43227);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_7 &&
	  wci_wciResponse_7$wget[33:32] == 2'd0 &&
	  !wci_respTimr_7_208_ULT_1_SL_wci_wTimeout_7_209_ETC___d5886 &&
	  wci_reqPend_7 == 2'd3)
	begin
	  v__h43316 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_7 &&
	  wci_wciResponse_7$wget[33:32] == 2'd0 &&
	  !wci_respTimr_7_208_ULT_1_SL_wci_wTimeout_7_209_ETC___d5886 &&
	  wci_reqPend_7 == 2'd3)
	$display("[%0d]: %m: WORKER CONTROL-OP   TIMEOUT", v__h43316);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_7 &&
	  wci_wciResponse_7$wget[33:32] == 2'd2 &&
	  wci_reqPend_7 == 2'd1)
	begin
	  v__h43540 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_7 &&
	  wci_wciResponse_7$wget[33:32] == 2'd2 &&
	  wci_reqPend_7 == 2'd1)
	$display("[%0d]: %m: WORKER CONFIG-WRITE RESPONSE-FAIL", v__h43540);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_7 &&
	  wci_wciResponse_7$wget[33:32] == 2'd2 &&
	  wci_reqPend_7 == 2'd2)
	begin
	  v__h43630 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_7 &&
	  wci_wciResponse_7$wget[33:32] == 2'd2 &&
	  wci_reqPend_7 == 2'd2)
	$display("[%0d]: %m: WORKER CONFIG-READ  RESPONSE-FAIL", v__h43630);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_7 &&
	  wci_wciResponse_7$wget[33:32] == 2'd2 &&
	  wci_reqPend_7 == 2'd3)
	begin
	  v__h43719 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_7 &&
	  wci_wciResponse_7$wget[33:32] == 2'd2 &&
	  wci_reqPend_7 == 2'd3)
	$display("[%0d]: %m: WORKER CONTROL-OP   RESPONSE-FAIL", v__h43719);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_7 &&
	  wci_wciResponse_7$wget[33:32] == 2'd3 &&
	  wci_reqPend_7 == 2'd1)
	begin
	  v__h43948 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_7 &&
	  wci_wciResponse_7$wget[33:32] == 2'd3 &&
	  wci_reqPend_7 == 2'd1)
	$display("[%0d]: %m: WORKER CONFIG-WRITE RESPONSE-ERR", v__h43948);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_7 &&
	  wci_wciResponse_7$wget[33:32] == 2'd3 &&
	  wci_reqPend_7 == 2'd2)
	begin
	  v__h44038 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_7 &&
	  wci_wciResponse_7$wget[33:32] == 2'd3 &&
	  wci_reqPend_7 == 2'd2)
	$display("[%0d]: %m: WORKER CONFIG-READ  RESPONSE-ERR", v__h44038);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_7 &&
	  wci_wciResponse_7$wget[33:32] == 2'd3 &&
	  wci_reqPend_7 == 2'd3)
	begin
	  v__h44127 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_7 &&
	  wci_wciResponse_7$wget[33:32] == 2'd3 &&
	  wci_reqPend_7 == 2'd3)
	$display("[%0d]: %m: WORKER CONTROL-OP   RESPONSE-ERR", v__h44127);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_8 &&
	  wci_wciResponse_8$wget[33:32] == 2'd0 &&
	  !wci_respTimr_8_348_ULT_1_SL_wci_wTimeout_8_349_ETC___d5887 &&
	  wci_reqPend_8 == 2'd1)
	begin
	  v__h47577 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_8 &&
	  wci_wciResponse_8$wget[33:32] == 2'd0 &&
	  !wci_respTimr_8_348_ULT_1_SL_wci_wTimeout_8_349_ETC___d5887 &&
	  wci_reqPend_8 == 2'd1)
	$display("[%0d]: %m: WORKER CONFIG-WRITE TIMEOUT", v__h47577);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_8 &&
	  wci_wciResponse_8$wget[33:32] == 2'd0 &&
	  !wci_respTimr_8_348_ULT_1_SL_wci_wTimeout_8_349_ETC___d5887 &&
	  wci_reqPend_8 == 2'd2)
	begin
	  v__h47667 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_8 &&
	  wci_wciResponse_8$wget[33:32] == 2'd0 &&
	  !wci_respTimr_8_348_ULT_1_SL_wci_wTimeout_8_349_ETC___d5887 &&
	  wci_reqPend_8 == 2'd2)
	$display("[%0d]: %m: WORKER CONFIG-READ  TIMEOUT", v__h47667);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_8 &&
	  wci_wciResponse_8$wget[33:32] == 2'd0 &&
	  !wci_respTimr_8_348_ULT_1_SL_wci_wTimeout_8_349_ETC___d5887 &&
	  wci_reqPend_8 == 2'd3)
	begin
	  v__h47756 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_8 &&
	  wci_wciResponse_8$wget[33:32] == 2'd0 &&
	  !wci_respTimr_8_348_ULT_1_SL_wci_wTimeout_8_349_ETC___d5887 &&
	  wci_reqPend_8 == 2'd3)
	$display("[%0d]: %m: WORKER CONTROL-OP   TIMEOUT", v__h47756);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_8 &&
	  wci_wciResponse_8$wget[33:32] == 2'd2 &&
	  wci_reqPend_8 == 2'd1)
	begin
	  v__h47980 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_8 &&
	  wci_wciResponse_8$wget[33:32] == 2'd2 &&
	  wci_reqPend_8 == 2'd1)
	$display("[%0d]: %m: WORKER CONFIG-WRITE RESPONSE-FAIL", v__h47980);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_8 &&
	  wci_wciResponse_8$wget[33:32] == 2'd2 &&
	  wci_reqPend_8 == 2'd2)
	begin
	  v__h48070 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_8 &&
	  wci_wciResponse_8$wget[33:32] == 2'd2 &&
	  wci_reqPend_8 == 2'd2)
	$display("[%0d]: %m: WORKER CONFIG-READ  RESPONSE-FAIL", v__h48070);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_8 &&
	  wci_wciResponse_8$wget[33:32] == 2'd2 &&
	  wci_reqPend_8 == 2'd3)
	begin
	  v__h48159 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_8 &&
	  wci_wciResponse_8$wget[33:32] == 2'd2 &&
	  wci_reqPend_8 == 2'd3)
	$display("[%0d]: %m: WORKER CONTROL-OP   RESPONSE-FAIL", v__h48159);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_8 &&
	  wci_wciResponse_8$wget[33:32] == 2'd3 &&
	  wci_reqPend_8 == 2'd1)
	begin
	  v__h48388 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_8 &&
	  wci_wciResponse_8$wget[33:32] == 2'd3 &&
	  wci_reqPend_8 == 2'd1)
	$display("[%0d]: %m: WORKER CONFIG-WRITE RESPONSE-ERR", v__h48388);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_8 &&
	  wci_wciResponse_8$wget[33:32] == 2'd3 &&
	  wci_reqPend_8 == 2'd2)
	begin
	  v__h48478 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_8 &&
	  wci_wciResponse_8$wget[33:32] == 2'd3 &&
	  wci_reqPend_8 == 2'd2)
	$display("[%0d]: %m: WORKER CONFIG-READ  RESPONSE-ERR", v__h48478);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_8 &&
	  wci_wciResponse_8$wget[33:32] == 2'd3 &&
	  wci_reqPend_8 == 2'd3)
	begin
	  v__h48567 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_8 &&
	  wci_wciResponse_8$wget[33:32] == 2'd3 &&
	  wci_reqPend_8 == 2'd3)
	$display("[%0d]: %m: WORKER CONTROL-OP   RESPONSE-ERR", v__h48567);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_9 &&
	  wci_wciResponse_9$wget[33:32] == 2'd0 &&
	  !wci_respTimr_9_488_ULT_1_SL_wci_wTimeout_9_489_ETC___d5888 &&
	  wci_reqPend_9 == 2'd1)
	begin
	  v__h52017 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_9 &&
	  wci_wciResponse_9$wget[33:32] == 2'd0 &&
	  !wci_respTimr_9_488_ULT_1_SL_wci_wTimeout_9_489_ETC___d5888 &&
	  wci_reqPend_9 == 2'd1)
	$display("[%0d]: %m: WORKER CONFIG-WRITE TIMEOUT", v__h52017);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_9 &&
	  wci_wciResponse_9$wget[33:32] == 2'd0 &&
	  !wci_respTimr_9_488_ULT_1_SL_wci_wTimeout_9_489_ETC___d5888 &&
	  wci_reqPend_9 == 2'd2)
	begin
	  v__h52107 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_9 &&
	  wci_wciResponse_9$wget[33:32] == 2'd0 &&
	  !wci_respTimr_9_488_ULT_1_SL_wci_wTimeout_9_489_ETC___d5888 &&
	  wci_reqPend_9 == 2'd2)
	$display("[%0d]: %m: WORKER CONFIG-READ  TIMEOUT", v__h52107);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_9 &&
	  wci_wciResponse_9$wget[33:32] == 2'd0 &&
	  !wci_respTimr_9_488_ULT_1_SL_wci_wTimeout_9_489_ETC___d5888 &&
	  wci_reqPend_9 == 2'd3)
	begin
	  v__h52196 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_9 &&
	  wci_wciResponse_9$wget[33:32] == 2'd0 &&
	  !wci_respTimr_9_488_ULT_1_SL_wci_wTimeout_9_489_ETC___d5888 &&
	  wci_reqPend_9 == 2'd3)
	$display("[%0d]: %m: WORKER CONTROL-OP   TIMEOUT", v__h52196);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_9 &&
	  wci_wciResponse_9$wget[33:32] == 2'd2 &&
	  wci_reqPend_9 == 2'd1)
	begin
	  v__h52420 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_9 &&
	  wci_wciResponse_9$wget[33:32] == 2'd2 &&
	  wci_reqPend_9 == 2'd1)
	$display("[%0d]: %m: WORKER CONFIG-WRITE RESPONSE-FAIL", v__h52420);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_9 &&
	  wci_wciResponse_9$wget[33:32] == 2'd2 &&
	  wci_reqPend_9 == 2'd2)
	begin
	  v__h52510 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_9 &&
	  wci_wciResponse_9$wget[33:32] == 2'd2 &&
	  wci_reqPend_9 == 2'd2)
	$display("[%0d]: %m: WORKER CONFIG-READ  RESPONSE-FAIL", v__h52510);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_9 &&
	  wci_wciResponse_9$wget[33:32] == 2'd2 &&
	  wci_reqPend_9 == 2'd3)
	begin
	  v__h52599 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_9 &&
	  wci_wciResponse_9$wget[33:32] == 2'd2 &&
	  wci_reqPend_9 == 2'd3)
	$display("[%0d]: %m: WORKER CONTROL-OP   RESPONSE-FAIL", v__h52599);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_9 &&
	  wci_wciResponse_9$wget[33:32] == 2'd3 &&
	  wci_reqPend_9 == 2'd1)
	begin
	  v__h52828 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_9 &&
	  wci_wciResponse_9$wget[33:32] == 2'd3 &&
	  wci_reqPend_9 == 2'd1)
	$display("[%0d]: %m: WORKER CONFIG-WRITE RESPONSE-ERR", v__h52828);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_9 &&
	  wci_wciResponse_9$wget[33:32] == 2'd3 &&
	  wci_reqPend_9 == 2'd2)
	begin
	  v__h52918 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_9 &&
	  wci_wciResponse_9$wget[33:32] == 2'd3 &&
	  wci_reqPend_9 == 2'd2)
	$display("[%0d]: %m: WORKER CONFIG-READ  RESPONSE-ERR", v__h52918);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_9 &&
	  wci_wciResponse_9$wget[33:32] == 2'd3 &&
	  wci_reqPend_9 == 2'd3)
	begin
	  v__h53007 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_9 &&
	  wci_wciResponse_9$wget[33:32] == 2'd3 &&
	  wci_reqPend_9 == 2'd3)
	$display("[%0d]: %m: WORKER CONTROL-OP   RESPONSE-ERR", v__h53007);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_10 &&
	  wci_wciResponse_10$wget[33:32] == 2'd0 &&
	  !wci_respTimr_10_628_ULT_1_SL_wci_wTimeout_10_6_ETC___d5889 &&
	  wci_reqPend_10 == 2'd1)
	begin
	  v__h56457 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_10 &&
	  wci_wciResponse_10$wget[33:32] == 2'd0 &&
	  !wci_respTimr_10_628_ULT_1_SL_wci_wTimeout_10_6_ETC___d5889 &&
	  wci_reqPend_10 == 2'd1)
	$display("[%0d]: %m: WORKER CONFIG-WRITE TIMEOUT", v__h56457);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_10 &&
	  wci_wciResponse_10$wget[33:32] == 2'd0 &&
	  !wci_respTimr_10_628_ULT_1_SL_wci_wTimeout_10_6_ETC___d5889 &&
	  wci_reqPend_10 == 2'd2)
	begin
	  v__h56547 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_10 &&
	  wci_wciResponse_10$wget[33:32] == 2'd0 &&
	  !wci_respTimr_10_628_ULT_1_SL_wci_wTimeout_10_6_ETC___d5889 &&
	  wci_reqPend_10 == 2'd2)
	$display("[%0d]: %m: WORKER CONFIG-READ  TIMEOUT", v__h56547);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_10 &&
	  wci_wciResponse_10$wget[33:32] == 2'd0 &&
	  !wci_respTimr_10_628_ULT_1_SL_wci_wTimeout_10_6_ETC___d5889 &&
	  wci_reqPend_10 == 2'd3)
	begin
	  v__h56636 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_10 &&
	  wci_wciResponse_10$wget[33:32] == 2'd0 &&
	  !wci_respTimr_10_628_ULT_1_SL_wci_wTimeout_10_6_ETC___d5889 &&
	  wci_reqPend_10 == 2'd3)
	$display("[%0d]: %m: WORKER CONTROL-OP   TIMEOUT", v__h56636);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_10 &&
	  wci_wciResponse_10$wget[33:32] == 2'd2 &&
	  wci_reqPend_10 == 2'd1)
	begin
	  v__h56860 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_10 &&
	  wci_wciResponse_10$wget[33:32] == 2'd2 &&
	  wci_reqPend_10 == 2'd1)
	$display("[%0d]: %m: WORKER CONFIG-WRITE RESPONSE-FAIL", v__h56860);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_10 &&
	  wci_wciResponse_10$wget[33:32] == 2'd2 &&
	  wci_reqPend_10 == 2'd2)
	begin
	  v__h56950 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_10 &&
	  wci_wciResponse_10$wget[33:32] == 2'd2 &&
	  wci_reqPend_10 == 2'd2)
	$display("[%0d]: %m: WORKER CONFIG-READ  RESPONSE-FAIL", v__h56950);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_10 &&
	  wci_wciResponse_10$wget[33:32] == 2'd2 &&
	  wci_reqPend_10 == 2'd3)
	begin
	  v__h57039 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_10 &&
	  wci_wciResponse_10$wget[33:32] == 2'd2 &&
	  wci_reqPend_10 == 2'd3)
	$display("[%0d]: %m: WORKER CONTROL-OP   RESPONSE-FAIL", v__h57039);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_10 &&
	  wci_wciResponse_10$wget[33:32] == 2'd3 &&
	  wci_reqPend_10 == 2'd1)
	begin
	  v__h57268 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_10 &&
	  wci_wciResponse_10$wget[33:32] == 2'd3 &&
	  wci_reqPend_10 == 2'd1)
	$display("[%0d]: %m: WORKER CONFIG-WRITE RESPONSE-ERR", v__h57268);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_10 &&
	  wci_wciResponse_10$wget[33:32] == 2'd3 &&
	  wci_reqPend_10 == 2'd2)
	begin
	  v__h57358 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_10 &&
	  wci_wciResponse_10$wget[33:32] == 2'd3 &&
	  wci_reqPend_10 == 2'd2)
	$display("[%0d]: %m: WORKER CONFIG-READ  RESPONSE-ERR", v__h57358);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_10 &&
	  wci_wciResponse_10$wget[33:32] == 2'd3 &&
	  wci_reqPend_10 == 2'd3)
	begin
	  v__h57447 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_10 &&
	  wci_wciResponse_10$wget[33:32] == 2'd3 &&
	  wci_reqPend_10 == 2'd3)
	$display("[%0d]: %m: WORKER CONTROL-OP   RESPONSE-ERR", v__h57447);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_11 &&
	  wci_wciResponse_11$wget[33:32] == 2'd0 &&
	  !wci_respTimr_11_768_ULT_1_SL_wci_wTimeout_11_7_ETC___d5890 &&
	  wci_reqPend_11 == 2'd1)
	begin
	  v__h60897 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_11 &&
	  wci_wciResponse_11$wget[33:32] == 2'd0 &&
	  !wci_respTimr_11_768_ULT_1_SL_wci_wTimeout_11_7_ETC___d5890 &&
	  wci_reqPend_11 == 2'd1)
	$display("[%0d]: %m: WORKER CONFIG-WRITE TIMEOUT", v__h60897);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_11 &&
	  wci_wciResponse_11$wget[33:32] == 2'd0 &&
	  !wci_respTimr_11_768_ULT_1_SL_wci_wTimeout_11_7_ETC___d5890 &&
	  wci_reqPend_11 == 2'd2)
	begin
	  v__h60987 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_11 &&
	  wci_wciResponse_11$wget[33:32] == 2'd0 &&
	  !wci_respTimr_11_768_ULT_1_SL_wci_wTimeout_11_7_ETC___d5890 &&
	  wci_reqPend_11 == 2'd2)
	$display("[%0d]: %m: WORKER CONFIG-READ  TIMEOUT", v__h60987);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_11 &&
	  wci_wciResponse_11$wget[33:32] == 2'd0 &&
	  !wci_respTimr_11_768_ULT_1_SL_wci_wTimeout_11_7_ETC___d5890 &&
	  wci_reqPend_11 == 2'd3)
	begin
	  v__h61076 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_11 &&
	  wci_wciResponse_11$wget[33:32] == 2'd0 &&
	  !wci_respTimr_11_768_ULT_1_SL_wci_wTimeout_11_7_ETC___d5890 &&
	  wci_reqPend_11 == 2'd3)
	$display("[%0d]: %m: WORKER CONTROL-OP   TIMEOUT", v__h61076);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_11 &&
	  wci_wciResponse_11$wget[33:32] == 2'd2 &&
	  wci_reqPend_11 == 2'd1)
	begin
	  v__h61300 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_11 &&
	  wci_wciResponse_11$wget[33:32] == 2'd2 &&
	  wci_reqPend_11 == 2'd1)
	$display("[%0d]: %m: WORKER CONFIG-WRITE RESPONSE-FAIL", v__h61300);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_11 &&
	  wci_wciResponse_11$wget[33:32] == 2'd2 &&
	  wci_reqPend_11 == 2'd2)
	begin
	  v__h61390 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_11 &&
	  wci_wciResponse_11$wget[33:32] == 2'd2 &&
	  wci_reqPend_11 == 2'd2)
	$display("[%0d]: %m: WORKER CONFIG-READ  RESPONSE-FAIL", v__h61390);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_11 &&
	  wci_wciResponse_11$wget[33:32] == 2'd2 &&
	  wci_reqPend_11 == 2'd3)
	begin
	  v__h61479 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_11 &&
	  wci_wciResponse_11$wget[33:32] == 2'd2 &&
	  wci_reqPend_11 == 2'd3)
	$display("[%0d]: %m: WORKER CONTROL-OP   RESPONSE-FAIL", v__h61479);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_11 &&
	  wci_wciResponse_11$wget[33:32] == 2'd3 &&
	  wci_reqPend_11 == 2'd1)
	begin
	  v__h61708 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_11 &&
	  wci_wciResponse_11$wget[33:32] == 2'd3 &&
	  wci_reqPend_11 == 2'd1)
	$display("[%0d]: %m: WORKER CONFIG-WRITE RESPONSE-ERR", v__h61708);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_11 &&
	  wci_wciResponse_11$wget[33:32] == 2'd3 &&
	  wci_reqPend_11 == 2'd2)
	begin
	  v__h61798 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_11 &&
	  wci_wciResponse_11$wget[33:32] == 2'd3 &&
	  wci_reqPend_11 == 2'd2)
	$display("[%0d]: %m: WORKER CONFIG-READ  RESPONSE-ERR", v__h61798);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_11 &&
	  wci_wciResponse_11$wget[33:32] == 2'd3 &&
	  wci_reqPend_11 == 2'd3)
	begin
	  v__h61887 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_11 &&
	  wci_wciResponse_11$wget[33:32] == 2'd3 &&
	  wci_reqPend_11 == 2'd3)
	$display("[%0d]: %m: WORKER CONTROL-OP   RESPONSE-ERR", v__h61887);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_12 &&
	  wci_wciResponse_12$wget[33:32] == 2'd0 &&
	  !wci_respTimr_12_908_ULT_1_SL_wci_wTimeout_12_9_ETC___d5891 &&
	  wci_reqPend_12 == 2'd1)
	begin
	  v__h65337 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_12 &&
	  wci_wciResponse_12$wget[33:32] == 2'd0 &&
	  !wci_respTimr_12_908_ULT_1_SL_wci_wTimeout_12_9_ETC___d5891 &&
	  wci_reqPend_12 == 2'd1)
	$display("[%0d]: %m: WORKER CONFIG-WRITE TIMEOUT", v__h65337);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_12 &&
	  wci_wciResponse_12$wget[33:32] == 2'd0 &&
	  !wci_respTimr_12_908_ULT_1_SL_wci_wTimeout_12_9_ETC___d5891 &&
	  wci_reqPend_12 == 2'd2)
	begin
	  v__h65427 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_12 &&
	  wci_wciResponse_12$wget[33:32] == 2'd0 &&
	  !wci_respTimr_12_908_ULT_1_SL_wci_wTimeout_12_9_ETC___d5891 &&
	  wci_reqPend_12 == 2'd2)
	$display("[%0d]: %m: WORKER CONFIG-READ  TIMEOUT", v__h65427);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_12 &&
	  wci_wciResponse_12$wget[33:32] == 2'd0 &&
	  !wci_respTimr_12_908_ULT_1_SL_wci_wTimeout_12_9_ETC___d5891 &&
	  wci_reqPend_12 == 2'd3)
	begin
	  v__h65516 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_12 &&
	  wci_wciResponse_12$wget[33:32] == 2'd0 &&
	  !wci_respTimr_12_908_ULT_1_SL_wci_wTimeout_12_9_ETC___d5891 &&
	  wci_reqPend_12 == 2'd3)
	$display("[%0d]: %m: WORKER CONTROL-OP   TIMEOUT", v__h65516);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_12 &&
	  wci_wciResponse_12$wget[33:32] == 2'd2 &&
	  wci_reqPend_12 == 2'd1)
	begin
	  v__h65740 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_12 &&
	  wci_wciResponse_12$wget[33:32] == 2'd2 &&
	  wci_reqPend_12 == 2'd1)
	$display("[%0d]: %m: WORKER CONFIG-WRITE RESPONSE-FAIL", v__h65740);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_12 &&
	  wci_wciResponse_12$wget[33:32] == 2'd2 &&
	  wci_reqPend_12 == 2'd2)
	begin
	  v__h65830 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_12 &&
	  wci_wciResponse_12$wget[33:32] == 2'd2 &&
	  wci_reqPend_12 == 2'd2)
	$display("[%0d]: %m: WORKER CONFIG-READ  RESPONSE-FAIL", v__h65830);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_12 &&
	  wci_wciResponse_12$wget[33:32] == 2'd2 &&
	  wci_reqPend_12 == 2'd3)
	begin
	  v__h65919 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_12 &&
	  wci_wciResponse_12$wget[33:32] == 2'd2 &&
	  wci_reqPend_12 == 2'd3)
	$display("[%0d]: %m: WORKER CONTROL-OP   RESPONSE-FAIL", v__h65919);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_12 &&
	  wci_wciResponse_12$wget[33:32] == 2'd3 &&
	  wci_reqPend_12 == 2'd1)
	begin
	  v__h66148 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_12 &&
	  wci_wciResponse_12$wget[33:32] == 2'd3 &&
	  wci_reqPend_12 == 2'd1)
	$display("[%0d]: %m: WORKER CONFIG-WRITE RESPONSE-ERR", v__h66148);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_12 &&
	  wci_wciResponse_12$wget[33:32] == 2'd3 &&
	  wci_reqPend_12 == 2'd2)
	begin
	  v__h66238 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_12 &&
	  wci_wciResponse_12$wget[33:32] == 2'd3 &&
	  wci_reqPend_12 == 2'd2)
	$display("[%0d]: %m: WORKER CONFIG-READ  RESPONSE-ERR", v__h66238);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_12 &&
	  wci_wciResponse_12$wget[33:32] == 2'd3 &&
	  wci_reqPend_12 == 2'd3)
	begin
	  v__h66327 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_12 &&
	  wci_wciResponse_12$wget[33:32] == 2'd3 &&
	  wci_reqPend_12 == 2'd3)
	$display("[%0d]: %m: WORKER CONTROL-OP   RESPONSE-ERR", v__h66327);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_13 &&
	  wci_wciResponse_13$wget[33:32] == 2'd0 &&
	  !wci_respTimr_13_048_ULT_1_SL_wci_wTimeout_13_0_ETC___d5892 &&
	  wci_reqPend_13 == 2'd1)
	begin
	  v__h69777 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_13 &&
	  wci_wciResponse_13$wget[33:32] == 2'd0 &&
	  !wci_respTimr_13_048_ULT_1_SL_wci_wTimeout_13_0_ETC___d5892 &&
	  wci_reqPend_13 == 2'd1)
	$display("[%0d]: %m: WORKER CONFIG-WRITE TIMEOUT", v__h69777);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_13 &&
	  wci_wciResponse_13$wget[33:32] == 2'd0 &&
	  !wci_respTimr_13_048_ULT_1_SL_wci_wTimeout_13_0_ETC___d5892 &&
	  wci_reqPend_13 == 2'd2)
	begin
	  v__h69867 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_13 &&
	  wci_wciResponse_13$wget[33:32] == 2'd0 &&
	  !wci_respTimr_13_048_ULT_1_SL_wci_wTimeout_13_0_ETC___d5892 &&
	  wci_reqPend_13 == 2'd2)
	$display("[%0d]: %m: WORKER CONFIG-READ  TIMEOUT", v__h69867);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_13 &&
	  wci_wciResponse_13$wget[33:32] == 2'd0 &&
	  !wci_respTimr_13_048_ULT_1_SL_wci_wTimeout_13_0_ETC___d5892 &&
	  wci_reqPend_13 == 2'd3)
	begin
	  v__h69956 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_13 &&
	  wci_wciResponse_13$wget[33:32] == 2'd0 &&
	  !wci_respTimr_13_048_ULT_1_SL_wci_wTimeout_13_0_ETC___d5892 &&
	  wci_reqPend_13 == 2'd3)
	$display("[%0d]: %m: WORKER CONTROL-OP   TIMEOUT", v__h69956);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_13 &&
	  wci_wciResponse_13$wget[33:32] == 2'd2 &&
	  wci_reqPend_13 == 2'd1)
	begin
	  v__h70180 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_13 &&
	  wci_wciResponse_13$wget[33:32] == 2'd2 &&
	  wci_reqPend_13 == 2'd1)
	$display("[%0d]: %m: WORKER CONFIG-WRITE RESPONSE-FAIL", v__h70180);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_13 &&
	  wci_wciResponse_13$wget[33:32] == 2'd2 &&
	  wci_reqPend_13 == 2'd2)
	begin
	  v__h70270 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_13 &&
	  wci_wciResponse_13$wget[33:32] == 2'd2 &&
	  wci_reqPend_13 == 2'd2)
	$display("[%0d]: %m: WORKER CONFIG-READ  RESPONSE-FAIL", v__h70270);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_13 &&
	  wci_wciResponse_13$wget[33:32] == 2'd2 &&
	  wci_reqPend_13 == 2'd3)
	begin
	  v__h70359 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_13 &&
	  wci_wciResponse_13$wget[33:32] == 2'd2 &&
	  wci_reqPend_13 == 2'd3)
	$display("[%0d]: %m: WORKER CONTROL-OP   RESPONSE-FAIL", v__h70359);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_13 &&
	  wci_wciResponse_13$wget[33:32] == 2'd3 &&
	  wci_reqPend_13 == 2'd1)
	begin
	  v__h70588 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_13 &&
	  wci_wciResponse_13$wget[33:32] == 2'd3 &&
	  wci_reqPend_13 == 2'd1)
	$display("[%0d]: %m: WORKER CONFIG-WRITE RESPONSE-ERR", v__h70588);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_13 &&
	  wci_wciResponse_13$wget[33:32] == 2'd3 &&
	  wci_reqPend_13 == 2'd2)
	begin
	  v__h70678 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_13 &&
	  wci_wciResponse_13$wget[33:32] == 2'd3 &&
	  wci_reqPend_13 == 2'd2)
	$display("[%0d]: %m: WORKER CONFIG-READ  RESPONSE-ERR", v__h70678);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_13 &&
	  wci_wciResponse_13$wget[33:32] == 2'd3 &&
	  wci_reqPend_13 == 2'd3)
	begin
	  v__h70767 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_13 &&
	  wci_wciResponse_13$wget[33:32] == 2'd3 &&
	  wci_reqPend_13 == 2'd3)
	$display("[%0d]: %m: WORKER CONTROL-OP   RESPONSE-ERR", v__h70767);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_14 &&
	  wci_wciResponse_14$wget[33:32] == 2'd0 &&
	  !wci_respTimr_14_188_ULT_1_SL_wci_wTimeout_14_1_ETC___d5893 &&
	  wci_reqPend_14 == 2'd1)
	begin
	  v__h74217 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_14 &&
	  wci_wciResponse_14$wget[33:32] == 2'd0 &&
	  !wci_respTimr_14_188_ULT_1_SL_wci_wTimeout_14_1_ETC___d5893 &&
	  wci_reqPend_14 == 2'd1)
	$display("[%0d]: %m: WORKER CONFIG-WRITE TIMEOUT", v__h74217);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_14 &&
	  wci_wciResponse_14$wget[33:32] == 2'd0 &&
	  !wci_respTimr_14_188_ULT_1_SL_wci_wTimeout_14_1_ETC___d5893 &&
	  wci_reqPend_14 == 2'd2)
	begin
	  v__h74307 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_14 &&
	  wci_wciResponse_14$wget[33:32] == 2'd0 &&
	  !wci_respTimr_14_188_ULT_1_SL_wci_wTimeout_14_1_ETC___d5893 &&
	  wci_reqPend_14 == 2'd2)
	$display("[%0d]: %m: WORKER CONFIG-READ  TIMEOUT", v__h74307);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_14 &&
	  wci_wciResponse_14$wget[33:32] == 2'd0 &&
	  !wci_respTimr_14_188_ULT_1_SL_wci_wTimeout_14_1_ETC___d5893 &&
	  wci_reqPend_14 == 2'd3)
	begin
	  v__h74396 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_14 &&
	  wci_wciResponse_14$wget[33:32] == 2'd0 &&
	  !wci_respTimr_14_188_ULT_1_SL_wci_wTimeout_14_1_ETC___d5893 &&
	  wci_reqPend_14 == 2'd3)
	$display("[%0d]: %m: WORKER CONTROL-OP   TIMEOUT", v__h74396);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_14 &&
	  wci_wciResponse_14$wget[33:32] == 2'd2 &&
	  wci_reqPend_14 == 2'd1)
	begin
	  v__h74620 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_14 &&
	  wci_wciResponse_14$wget[33:32] == 2'd2 &&
	  wci_reqPend_14 == 2'd1)
	$display("[%0d]: %m: WORKER CONFIG-WRITE RESPONSE-FAIL", v__h74620);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_14 &&
	  wci_wciResponse_14$wget[33:32] == 2'd2 &&
	  wci_reqPend_14 == 2'd2)
	begin
	  v__h74710 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_14 &&
	  wci_wciResponse_14$wget[33:32] == 2'd2 &&
	  wci_reqPend_14 == 2'd2)
	$display("[%0d]: %m: WORKER CONFIG-READ  RESPONSE-FAIL", v__h74710);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_14 &&
	  wci_wciResponse_14$wget[33:32] == 2'd2 &&
	  wci_reqPend_14 == 2'd3)
	begin
	  v__h74799 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_14 &&
	  wci_wciResponse_14$wget[33:32] == 2'd2 &&
	  wci_reqPend_14 == 2'd3)
	$display("[%0d]: %m: WORKER CONTROL-OP   RESPONSE-FAIL", v__h74799);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_14 &&
	  wci_wciResponse_14$wget[33:32] == 2'd3 &&
	  wci_reqPend_14 == 2'd1)
	begin
	  v__h75028 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_14 &&
	  wci_wciResponse_14$wget[33:32] == 2'd3 &&
	  wci_reqPend_14 == 2'd1)
	$display("[%0d]: %m: WORKER CONFIG-WRITE RESPONSE-ERR", v__h75028);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_14 &&
	  wci_wciResponse_14$wget[33:32] == 2'd3 &&
	  wci_reqPend_14 == 2'd2)
	begin
	  v__h75118 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_14 &&
	  wci_wciResponse_14$wget[33:32] == 2'd3 &&
	  wci_reqPend_14 == 2'd2)
	$display("[%0d]: %m: WORKER CONFIG-READ  RESPONSE-ERR", v__h75118);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_14 &&
	  wci_wciResponse_14$wget[33:32] == 2'd3 &&
	  wci_reqPend_14 == 2'd3)
	begin
	  v__h75207 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wci_wrkBusy_14 &&
	  wci_wciResponse_14$wget[33:32] == 2'd3 &&
	  wci_reqPend_14 == 2'd3)
	$display("[%0d]: %m: WORKER CONTROL-OP   RESPONSE-ERR", v__h75207);
  end
  // synopsys translate_on
endmodule  // mkOCCP

