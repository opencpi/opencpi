-- THIS FILE WAS ORIGINALLY GENERATED ON Mon Oct  1 17:09:18 2012 EDT
-- BASED ON THE FILE: gen/fsk_mod_complex.xml
-- YOU *ARE* EXPECTED TO EDIT IT
-- This file initially contains the architecture skeleton for worker: fsk_mod_complex

library IEEE; use IEEE.std_logic_1164.all; use ieee.numeric_std.all;
library ocpi; use ocpi.types.all; -- remove this to avoid all ocpi name collisions
architecture rtl of fsk_mod_complex_worker is
begin
end rtl;
