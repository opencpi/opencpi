// THIS FILE WAS ORIGINALLY GENERATED ON Thu Sep 20 16:14:53 2012 EDT
// BASED ON THE FILE: sym_fir_real.xml
// YOU ARE EXPECTED TO EDIT IT
// This file contains the implementation skeleton for worker: sym_fir_real

`include "sym_fir_real-impl.vh"



endmodule //sym_fir_real
