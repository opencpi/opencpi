(* box_type="user_black_box" *)
module mkUUID(uuid);
  // value method uuid
  output [511 : 0] uuid;
endmodule  // mkUUID

