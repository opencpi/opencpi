// THIS FILE WAS ORIGINALLY GENERATED ON Thu Sep 20 16:14:52 2012 EDT
// BASED ON THE FILE: cic_lpfilter_complex.xml
// YOU ARE EXPECTED TO EDIT IT
// This file contains the implementation skeleton for worker: cic_lpfilter_complex

`include "cic_lpfilter_complex-impl.vh"



endmodule //cic_lpfilter_complex
