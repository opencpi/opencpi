../../../optical_flow_pyr_lk.rcc/target-linux-c6-x86_64/generics.vhd