../../../../assets/hdl/devices/ad9361_spi.hdl/signals.vhd