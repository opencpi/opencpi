-- THIS FILE WAS ORIGINALLY GENERATED ON Tue Apr 16 15:06:04 2013 EDT
-- BASED ON THE FILE: capture_vhdl.xml
-- YOU *ARE* EXPECTED TO EDIT IT
-- This file initially contains the architecture skeleton for worker: capture_vhdl

library IEEE; use IEEE.std_logic_1164.all; use ieee.numeric_std.all;
library ocpi; use ocpi.types.all; -- remove this to avoid all ocpi name collisions
architecture rtl of capture_vhdl_worker is
begin
end rtl;
