-- This file is protected by Copyright. Please refer to the COPYRIGHT file
-- distributed with this source distribution.
--
-- This file is part of OpenCPI <http:--www.opencpi.org>
--
-- OpenCPI is free software: you can redistribute it and/or modify it under the
-- terms of the GNU Lesser General Public License as published by the Free
-- Software Foundation, either version 3 of the License, or (at your option) any
-- later version.
--
-- OpenCPI is distributed in the hope that it will be useful, but WITHOUT ANY
-- WARRANTY; without even the implied warranty of MERCHANTABILITY or FITNESS FOR
-- A PARTICULAR PURPOSE. See the GNU Lesser General Public License for more
-- details.
--
-- You should have received a copy of the GNU Lesser General Public License
-- along with this program. If not, see <http:--www.gnu.org/licenses/>.

-- This file is our wrapper around the processing_system8 IP as generated by
-- ps8.tcl.
-- There is no logic here, just providing a simpler interface for the platform worker
-- that uses it.
library IEEE; use IEEE.std_logic_1164.all; use ieee.numeric_std.all;
library ocpi; use ocpi.types.all; -- remove this to avoid all ocpi name collisions
library zynq_ultra; use zynq_ultra.zynq_ultra_pkg.all;
library axi; use axi.axi_pkg.all;
library zynq_ultra; use zynq_ultra.zynq_ultra_ps_e_wrap.all;
entity zynq_ultra_ps_e is
  port(
    ps_in        : in    pl2ps_t;
    ps_out       : out   ps2pl_t;
    m_axi_hp_in  : in    m_axi_hp_in_array_t(0 to C_M_AXI_HP_COUNT-1);
    m_axi_hp_out : out   m_axi_hp_out_array_t(0 to C_M_AXI_HP_COUNT-1);
    s_axi_hp_in  : in    s_axi_hp_in_array_t(0 to C_S_AXI_HP_COUNT-1);
    s_axi_hp_out : out   s_axi_hp_out_array_t(0 to C_S_AXI_HP_COUNT-1)
    );
end entity zynq_ultra_ps_e;
architecture rtl of zynq_ultra_ps_e is
  -- Various SLV arrays of different SLV widths for use below
  type vec_49_array_t is array (natural range <>) of std_logic_vector(48 downto 0);
  type vec_40_array_t is array (natural range <>) of std_logic_vector(39 downto 0);
  type vec_32_array_t is array (natural range <>) of std_logic_vector(31 downto 0);
  type vec_16_array_t is array (natural range <>) of std_logic_vector(15 downto 0);
  type vec_8_array_t is array (natural range <>) of std_logic_vector(7 downto 0);
  type vec_6_array_t is array (natural range <>) of std_logic_vector(5 downto 0);
  type vec_4_array_t is array (natural range <>) of std_logic_vector(3 downto 0);

  -- Some AXI signals have bit-width mismatches between the UltraScale PS8 and
  -- the OpenCPI AXI primitive. These intermediate signals below are used to
  -- compensate for the mismatches by leaving higher-order unused signals open
  -- or tied to '0'
  signal maxigp_awaddrs : vec_40_array_t(0 to C_M_AXI_HP_COUNT-1);
  signal maxigp_awlens  : vec_8_array_t (0 to C_M_AXI_HP_COUNT-1);
  signal maxigp_awids   : vec_16_array_t(0 to C_M_AXI_HP_COUNT-1);

  signal maxigp_araddrs : vec_40_array_t(0 to C_M_AXI_HP_COUNT-1);
  signal maxigp_arlens  : vec_8_array_t (0 to C_M_AXI_HP_COUNT-1);
  signal maxigp_arids   : vec_16_array_t(0 to C_M_AXI_HP_COUNT-1);

  signal maxigp_bids    : vec_16_array_t(0 to C_M_AXI_HP_COUNT-1);
  signal maxigp_rids    : vec_16_array_t(0 to C_M_AXI_HP_COUNT-1);

  signal saxigp_awaddrs : vec_49_array_t(0 to C_S_AXI_HP_COUNT-1);
  signal saxigp_awlens  : vec_8_array_t (0 to C_S_AXI_HP_COUNT-1);

  signal saxigp_araddrs : vec_49_array_t(0 to C_S_AXI_HP_COUNT-1);
  signal saxigp_arlens  : vec_8_array_t (0 to C_S_AXI_HP_COUNT-1);

begin

  -- The generate blocks below adapt bit-widths for the 40-bit address space
  -- of the ZynqMP's AXI to the 32-bit address space of the OpenCPI AXI primitive
  -- (tie higher-order unused signals to '0' and connect only needed ones)
  m : for i in 0 to C_M_AXI_HP_COUNT-1 generate
    m_axi_hp_out(i).ARESETN <= '1';
    m_axi_hp_out(i).W.ID <= (others => '0');

    m_axi_hp_out(i).AW.ADDR <= maxigp_awaddrs(i)(31 downto 0);
    m_axi_hp_out(i).AW.LEN <= maxigp_awlens(i)(3 downto 0);
    m_axi_hp_out(i).AW.ID <= maxigp_awids(i)(11 downto 0);
    m_axi_hp_out(i).AW.LOCK(1) <= '0';
    m_axi_hp_out(i).AW.ISSUECAP1_EN <= '0';
    m_axi_hp_out(i).AW.COUNT <= (others => '0');

    m_axi_hp_out(i).AR.ADDR <= maxigp_araddrs(i)(31 downto 0);
    m_axi_hp_out(i).AR.LEN <= maxigp_arlens(i)(3 downto 0);
    m_axi_hp_out(i).AR.ID <= maxigp_arids(i)(11 downto 0);
    m_axi_hp_out(i).AR.ISSUECAP1_EN <= '0';
    m_axi_hp_out(i).AR.COUNT <= (others => '0');

    maxigp_bids(i)(11 downto 0)  <= m_axi_hp_in(0).B.ID;
    maxigp_bids(i)(15 downto 12) <= (others =>'0');

    maxigp_rids(i)(11 downto 0) <= m_axi_hp_in(0).R.ID;
    maxigp_rids(i)(15 downto 12) <= (others =>'0');
  end generate;

  s : for i in 0 to C_S_AXI_HP_COUNT-1 generate
    s_axi_hp_out(i).ARESETN <= '1';

    saxigp_awaddrs(i)(31 downto 0)  <= s_axi_hp_in(0).AW.ADDR;
    saxigp_awaddrs(i)(48 downto 32) <= (others =>'0');
    saxigp_awlens(i)(3 downto 0)  <= s_axi_hp_in(0).AW.LEN;
    saxigp_awlens(i)(7 downto 4) <= (others =>'0');
    s_axi_hp_out(i).AW.COUNT <= (others => '0');

    saxigp_araddrs(i)(31 downto 0)  <= s_axi_hp_in(0).AR.ADDR;
    saxigp_araddrs(i)(48 downto 32) <= (others =>'0');
    saxigp_arlens(i)(3 downto 0)  <= s_axi_hp_in(0).AR.LEN;
    saxigp_arlens(i)(7 downto 4) <= (others =>'0');
    s_axi_hp_out(i).AR.COUNT <= (others => '0');

  end generate;

  -- Connect the Verilog PS8 wrapper to the VHDL axi records to abstract the interface
  ps : zynq_ultra_ps_e_0
    port map(
-- maxigp0
      maxihpm0_fpd_aclk => m_axi_hp_in(0).ACLK,
      maxigp0_awid => maxigp_awids(0), --[15:0]
      maxigp0_awaddr => maxigp_awaddrs(0), --[39:0]
      maxigp0_awlen => maxigp_awlens(0), --[7:0]
      maxigp0_awsize => m_axi_hp_out(0).AW.SIZE, --[2:0]
      maxigp0_awburst => m_axi_hp_out(0).AW.BURST, --[1:0]
      maxigp0_awlock => m_axi_hp_out(0).AW.LOCK(0),
      maxigp0_awcache => m_axi_hp_out(0).AW.CACHE, --[3:0]
      maxigp0_awprot => m_axi_hp_out(0).AW.PROT, --[2:0]
      maxigp0_awvalid => m_axi_hp_out(0).AW.VALID,
      maxigp0_awuser => open, --[15:0]
      maxigp0_awready => m_axi_hp_in(0).AW.READY,
      maxigp0_wdata => m_axi_hp_out(0).W.DATA, --[C_MAXIGP0_DATA_WIDTH-1 :0]
      maxigp0_wstrb => m_axi_hp_out(0).W.STRB, --[(C_MAXIGP0_DATA_WIDTH/8)-1 :0]
      maxigp0_wlast => m_axi_hp_out(0).W.LAST,
      maxigp0_wvalid => m_axi_hp_out(0).W.VALID,
      maxigp0_wready => m_axi_hp_in(0).W.READY,
      maxigp0_bid => maxigp_bids(0), --[15:0]
      maxigp0_bresp => m_axi_hp_in(0).B.RESP, --[1:0]
      maxigp0_bvalid => m_axi_hp_in(0).B.VALID,
      maxigp0_bready => m_axi_hp_out(0).B.READY,
      maxigp0_arid => maxigp_arids(0), --[15:0]
      maxigp0_araddr => maxigp_araddrs(0), --[39:0]
      maxigp0_arlen => maxigp_arlens(0), --[7:0]
      maxigp0_arsize => m_axi_hp_out(0).AR.SIZE, --[2:0]
      maxigp0_arburst => m_axi_hp_out(0).AR.BURST, --[1:0]
      maxigp0_arlock => m_axi_hp_out(0).AR.LOCK(0),
      maxigp0_arcache => m_axi_hp_out(0).AR.CACHE, --[3:0]
      maxigp0_arprot => m_axi_hp_out(0).AR.PROT, --[2:0]
      maxigp0_arvalid => m_axi_hp_out(0).AR.VALID,
      maxigp0_aruser => open, --[15:0]
      maxigp0_arready => m_axi_hp_in(0).AR.READY,
      maxigp0_rid => maxigp_rids(0), --[15:0]
      maxigp0_rdata => m_axi_hp_in(0).R.DATA, --[C_MAXIGP0_DATA_WIDTH-1 :0]
      maxigp0_rresp => m_axi_hp_in(0).R.RESP, --[1:0]
      maxigp0_rlast => m_axi_hp_in(0).R.LAST,
      maxigp0_rvalid => m_axi_hp_in(0).R.VALID,
      maxigp0_rready => m_axi_hp_out(0).R.READY,
      maxigp0_awqos => m_axi_hp_out(0).AW.QOS, --[3:0]
      maxigp0_arqos => m_axi_hp_out(0).AR.QOS, --[3:0]

-- maxigp1
      maxihpm1_fpd_aclk => m_axi_hp_in(1).ACLK,
      maxigp1_awid => maxigp_awids(1),
      maxigp1_awaddr => maxigp_awaddrs(1),
      maxigp1_awlen => maxigp_awlens(1),
      maxigp1_awsize => m_axi_hp_out(1).AW.SIZE, --[2:0]
      maxigp1_awburst => m_axi_hp_out(1).AW.BURST, --[1:0]
      maxigp1_awlock => m_axi_hp_out(1).AW.LOCK(0),
      maxigp1_awcache => m_axi_hp_out(1).AW.CACHE, --[3:0]
      maxigp1_awprot => m_axi_hp_out(1).AW.PROT, --[2:0]
      maxigp1_awvalid => m_axi_hp_out(1).AW.VALID,
      maxigp1_awuser => open, --[15:0]
      maxigp1_awready => m_axi_hp_in(1).AW.READY,
      maxigp1_wdata => m_axi_hp_out(1).W.DATA, --[C_MAXIGP1_DATA_WIDTH-1 :0]
      maxigp1_wstrb => m_axi_hp_out(1).W.STRB, --[(C_MAXIGP1_DATA_WIDTH/8)-1 :0]
      maxigp1_wlast => m_axi_hp_out(1).W.LAST,
      maxigp1_wvalid => m_axi_hp_out(1).W.VALID,
      maxigp1_wready => m_axi_hp_in(1).W.READY,
      maxigp1_bid => maxigp_bids(1), --m_axi_hp_in(1).B.ID, --[15:0]
      maxigp1_bresp => m_axi_hp_in(1).B.RESP, --[1:0]
      maxigp1_bvalid => m_axi_hp_in(1).B.VALID,
      maxigp1_bready => m_axi_hp_out(1).B.READY,
      maxigp1_arid => maxigp_arids(1),
      maxigp1_araddr => maxigp_araddrs(1),
      maxigp1_arlen => maxigp_arlens(1),
      maxigp1_arsize => m_axi_hp_out(1).AR.SIZE, --[2:0]
      maxigp1_arburst => m_axi_hp_out(1).AR.BURST, --[1:0]
      maxigp1_arlock => m_axi_hp_out(1).AR.LOCK(0),
      maxigp1_arprot => m_axi_hp_out(1).AR.PROT, --[2:0]
      maxigp1_arcache => m_axi_hp_out(1).AR.CACHE, --[3:0]
      maxigp1_arvalid => m_axi_hp_out(1).AR.VALID,
      maxigp1_aruser => open, --[15:0]
      maxigp1_arready => m_axi_hp_in(1).AR.READY,
      maxigp1_rid => maxigp_rids(1), --[15:0]
      maxigp1_rdata => m_axi_hp_in(1).R.DATA, --[C_MAXIGP1_DATA_WIDTH-1 :0]
      maxigp1_rresp => m_axi_hp_in(1).R.RESP, --[1:0]
      maxigp1_rlast => m_axi_hp_in(1).R.LAST,
      maxigp1_rvalid => m_axi_hp_in(1).R.VALID,
      maxigp1_rready => m_axi_hp_out(1).R.READY,
      maxigp1_awqos => m_axi_hp_out(1).AW.QOS, --[3:0]
      maxigp1_arqos => m_axi_hp_out(1).AR.QOS, --[3:0]
-- saxigp2
      saxihp0_fpd_aclk => s_axi_hp_in(0).ACLK,
      saxigp2_aruser => '0',
      saxigp2_awuser => '0',
      saxigp2_awid => s_axi_hp_in(0).AW.ID(5 downto 0), --[5:0]
      saxigp2_awaddr => saxigp_awaddrs(0), --[48:0]
      saxigp2_awlen => saxigp_awlens(0), --[7:0]
      saxigp2_awsize => s_axi_hp_in(0).AW.SIZE, --[2:0]
      saxigp2_awburst => s_axi_hp_in(0).AW.BURST, --[1:0]
      saxigp2_awlock => s_axi_hp_in(0).AW.LOCK(0),
      saxigp2_awcache => s_axi_hp_in(0).AW.CACHE, --[3:0]
      saxigp2_awprot => s_axi_hp_in(0).AW.PROT, --[2:0]
      saxigp2_awvalid => s_axi_hp_in(0).AW.VALID,
      saxigp2_awready => s_axi_hp_out(0).AW.READY,
      saxigp2_wdata => s_axi_hp_in(0).W.DATA, --[C_SAXIGP2_DATA_WIDTH-1:0]
      saxigp2_wstrb => s_axi_hp_in(0).W.STRB, --[(C_SAXIGP2_DATA_WIDTH/8) -1 :0]
      saxigp2_wlast => s_axi_hp_in(0).W.LAST,
      saxigp2_wvalid => s_axi_hp_in(0).W.VALID,
      saxigp2_wready => s_axi_hp_out(0).W.READY,
      saxigp2_bid => s_axi_hp_out(0).B.ID(5 downto 0), --[5:0]
      saxigp2_bresp => s_axi_hp_out(0).B.RESP, --[1:0]
      saxigp2_bvalid => s_axi_hp_out(0).B.VALID,
      saxigp2_bready => s_axi_hp_in(0).B.READY,
      saxigp2_arid => s_axi_hp_in(0).AR.ID(5 downto 0), --[5:0]
      saxigp2_araddr => saxigp_araddrs(0), --[48:0]
      saxigp2_arlen => saxigp_arlens(0), --[7:0]
      saxigp2_arsize => s_axi_hp_in(0).AR.SIZE, --[2:0]
      saxigp2_arburst => s_axi_hp_in(0).AR.BURST, --[1:0]
      saxigp2_arlock => s_axi_hp_in(0).AR.LOCK(0),
      saxigp2_arcache => s_axi_hp_in(0).AR.CACHE, --[3:0]
      saxigp2_arprot => s_axi_hp_in(0).AR.PROT, --[2:0]
      saxigp2_arvalid => s_axi_hp_in(0).AR.VALID,
      saxigp2_arready => s_axi_hp_out(0).AR.READY,
      saxigp2_rid => s_axi_hp_out(0).R.ID(5 downto 0), --[5:0]
      saxigp2_rdata => s_axi_hp_out(0).R.DATA, --[C_SAXIGP2_DATA_WIDTH-1:0]
      saxigp2_rresp => s_axi_hp_out(0).R.RESP, --[1:0]
      saxigp2_rlast => s_axi_hp_out(0).R.LAST,
      saxigp2_rvalid => s_axi_hp_out(0).R.VALID,
      saxigp2_rready => s_axi_hp_in(0).R.READY,
      saxigp2_awqos => s_axi_hp_in(0).AW.QOS, --[3:0]
      saxigp2_arqos => s_axi_hp_in(0).AR.QOS, --[3:0]
-- saxigp3
      saxihp1_fpd_aclk => s_axi_hp_in(1).ACLK,
      saxigp3_aruser => '0',
      saxigp3_awuser => '0',
      saxigp3_awid => s_axi_hp_in(1).AW.ID(5 downto 0), --[5:0]
      saxigp3_awaddr => saxigp_awaddrs(1), --[48:0]
      saxigp3_awlen => saxigp_awlens(1), --[7:0]
      saxigp3_awsize => s_axi_hp_in(1).AW.SIZE, --[2:0]
      saxigp3_awburst => s_axi_hp_in(1).AW.BURST, --[1:0]
      saxigp3_awlock => s_axi_hp_in(1).AW.LOCK(0),
      saxigp3_awcache => s_axi_hp_in(1).AW.CACHE, --[3:0]
      saxigp3_awprot => s_axi_hp_in(1).AW.PROT, --[2:0]
      saxigp3_awvalid => s_axi_hp_in(1).AW.VALID,
      saxigp3_awready => s_axi_hp_out(1).AW.READY,
      saxigp3_wdata => s_axi_hp_in(1).W.DATA, --[C_SAXIGP3_DATA_WIDTH-1:0]
      saxigp3_wstrb => s_axi_hp_in(1).W.STRB, --[(C_SAXIGP3_DATA_WIDTH/8) -1 :0]
      saxigp3_wlast => s_axi_hp_in(1).W.LAST,
      saxigp3_wvalid => s_axi_hp_in(1).W.VALID,
      saxigp3_wready => s_axi_hp_out(1).W.READY,
      saxigp3_bid => s_axi_hp_out(1).B.ID(5 downto 0), --[5:0]
      saxigp3_bresp => s_axi_hp_out(1).B.RESP, --[1:0]
      saxigp3_bvalid => s_axi_hp_out(1).B.VALID,
      saxigp3_bready => s_axi_hp_in(1).B.READY,
      saxigp3_arid => s_axi_hp_in(1).AR.ID(5 downto 0), --[5:0]
      saxigp3_araddr => saxigp_araddrs(1), --[48:0]
      saxigp3_arlen => saxigp_arlens(1), --[7:0]
      saxigp3_arsize => s_axi_hp_in(1).AR.SIZE, --[2:0]
      saxigp3_arburst => s_axi_hp_in(1).AR.BURST, --[1:0]
      saxigp3_arlock => s_axi_hp_in(1).AR.LOCK(0),
      saxigp3_arcache => s_axi_hp_in(1).AR.CACHE, --[3:0]
      saxigp3_arprot => s_axi_hp_in(1).AR.PROT, --[2:0]
      saxigp3_arvalid => s_axi_hp_in(1).AR.VALID,
      saxigp3_arready => s_axi_hp_out(1).AR.READY,
      saxigp3_rid => s_axi_hp_out(1).R.ID(5 downto 0), --[5:0]
      saxigp3_rdata => s_axi_hp_out(1).R.DATA, --[C_SAXIGP3_DATA_WIDTH-1:0]
      saxigp3_rresp => s_axi_hp_out(1).R.RESP, --[1:0]
      saxigp3_rlast => s_axi_hp_out(1).R.LAST,
      saxigp3_rvalid => s_axi_hp_out(1).R.VALID,
      saxigp3_rready => s_axi_hp_in(1).R.READY,
      saxigp3_awqos => s_axi_hp_in(1).AW.QOS, --[3:0]
      saxigp3_arqos => s_axi_hp_in(1).AR.QOS, --[3:0]
-- saxigp4
      saxihp2_fpd_aclk => s_axi_hp_in(2).ACLK,
      saxigp4_aruser => '0',
      saxigp4_awuser => '0',
      saxigp4_awid => s_axi_hp_in(2).AW.ID(5 downto 0), --[5:0]
      saxigp4_awaddr => saxigp_awaddrs(2), --[48:0]
      saxigp4_awlen => saxigp_awlens(2), --[7:0]
      saxigp4_awsize => s_axi_hp_in(2).AW.SIZE, --[2:0]
      saxigp4_awburst => s_axi_hp_in(2).AW.BURST, --[1:0]
      saxigp4_awlock => s_axi_hp_in(2).AW.LOCK(0),
      saxigp4_awcache => s_axi_hp_in(2).AW.CACHE, --[3:0]
      saxigp4_awprot => s_axi_hp_in(2).AW.PROT, --[2:0]
      saxigp4_awvalid => s_axi_hp_in(2).AW.VALID,
      saxigp4_awready => s_axi_hp_out(2).AW.READY,
      saxigp4_wdata => s_axi_hp_in(2).W.DATA, --[C_SAXIGP4_DATA_WIDTH-1:0]
      saxigp4_wstrb => s_axi_hp_in(2).W.STRB, --[(C_SAXIGP4_DATA_WIDTH/8) -1 :0]
      saxigp4_wlast => s_axi_hp_in(2).W.LAST,
      saxigp4_wvalid => s_axi_hp_in(2).W.VALID,
      saxigp4_wready => s_axi_hp_out(2).W.READY,
      saxigp4_bid => s_axi_hp_out(2).B.ID(5 downto 0), --[5:0]
      saxigp4_bresp => s_axi_hp_out(2).B.RESP, --[1:0]
      saxigp4_bvalid => s_axi_hp_out(2).B.VALID,
      saxigp4_bready => s_axi_hp_in(2).B.READY,
      saxigp4_arid => s_axi_hp_in(2).AR.ID(5 downto 0), --[5:0]
      saxigp4_araddr => saxigp_araddrs(2), --[48:0]
      saxigp4_arlen => saxigp_arlens(2), --[7:0]
      saxigp4_arsize => s_axi_hp_in(2).AR.SIZE, --[2:0]
      saxigp4_arburst => s_axi_hp_in(2).AR.BURST, --[1:0]
      saxigp4_arlock => s_axi_hp_in(2).AR.LOCK(0),
      saxigp4_arcache => s_axi_hp_in(2).AR.CACHE, --[3:0]
      saxigp4_arprot => s_axi_hp_in(2).AR.PROT, --[2:0]
      saxigp4_arvalid => s_axi_hp_in(2).AR.VALID,
      saxigp4_arready => s_axi_hp_out(2).AR.READY,
      saxigp4_rid => s_axi_hp_out(2).R.ID(5 downto 0), --[5:0]
      saxigp4_rdata => s_axi_hp_out(2).R.DATA, --[C_SAXIGP4_DATA_WIDTH-1:0]
      saxigp4_rresp => s_axi_hp_out(2).R.RESP, --[1:0]
      saxigp4_rlast => s_axi_hp_out(2).R.LAST,
      saxigp4_rvalid => s_axi_hp_out(2).R.VALID,
      saxigp4_rready => s_axi_hp_in(2).R.READY,
      saxigp4_awqos => s_axi_hp_in(2).AW.QOS, --[3:0]
      saxigp4_arqos => s_axi_hp_in(2).AR.QOS, --[3:0]
-- saxigp5
      saxihp3_fpd_aclk => s_axi_hp_in(3).ACLK,
      saxigp5_aruser => '0',
      saxigp5_awuser => '0',
      saxigp5_awid => s_axi_hp_in(3).AW.ID(5 downto 0), --[5:0]
      saxigp5_awaddr => saxigp_awaddrs(3), --[48:0]
      saxigp5_awlen => saxigp_awlens(3), --[7:0]
      saxigp5_awsize => s_axi_hp_in(3).AW.SIZE, --[2:0]
      saxigp5_awburst => s_axi_hp_in(3).AW.BURST, --[1:0]
      saxigp5_awlock => s_axi_hp_in(3).AW.LOCK(0),
      saxigp5_awcache => s_axi_hp_in(3).AW.CACHE, --[3:0]
      saxigp5_awprot => s_axi_hp_in(3).AW.PROT, --[2:0]
      saxigp5_awvalid => s_axi_hp_in(3).AW.VALID,
      saxigp5_awready => s_axi_hp_out(3).AW.READY,
      saxigp5_wdata => s_axi_hp_in(3).W.DATA, --[C_SAXIGP5_DATA_WIDTH-1:0]
      saxigp5_wstrb => s_axi_hp_in(3).W.STRB, --[(C_SAXIGP5_DATA_WIDTH/8) -1 :0]
      saxigp5_wlast => s_axi_hp_in(3).W.LAST,
      saxigp5_wvalid => s_axi_hp_in(3).W.VALID,
      saxigp5_wready => s_axi_hp_out(3).W.READY,
      saxigp5_bid => s_axi_hp_out(3).B.ID(5 downto 0), --[5:0]
      saxigp5_bresp => s_axi_hp_out(3).B.RESP, --[1:0]
      saxigp5_bvalid => s_axi_hp_out(3).B.VALID,
      saxigp5_bready => s_axi_hp_in(3).B.READY,
      saxigp5_arid => s_axi_hp_in(3).AR.ID(5 downto 0), --[5:0]
      saxigp5_araddr => saxigp_araddrs(3), --[48:0]
      saxigp5_arlen => saxigp_arlens(3), --[7:0]
      saxigp5_arsize => s_axi_hp_in(3).AR.SIZE, --[2:0]
      saxigp5_arburst => s_axi_hp_in(3).AR.BURST, --[1:0]
      saxigp5_arlock => s_axi_hp_in(3).AR.LOCK(0),
      saxigp5_arcache => s_axi_hp_in(3).AR.CACHE, --[3:0]
      saxigp5_arprot => s_axi_hp_in(3).AR.PROT, --[2:0]
      saxigp5_arvalid => s_axi_hp_in(3).AR.VALID,
      saxigp5_arready => s_axi_hp_out(3).AR.READY,
      saxigp5_rid => s_axi_hp_out(3).R.ID(5 downto 0), --[5:0]
      saxigp5_rdata => s_axi_hp_out(3).R.DATA, --[C_SAXIGP5_DATA_WIDTH-1:0]
      saxigp5_rresp => s_axi_hp_out(3).R.RESP, --[1:0]
      saxigp5_rlast => s_axi_hp_out(3).R.LAST,
      saxigp5_rvalid => s_axi_hp_out(3).R.VALID,
      saxigp5_rready => s_axi_hp_in(3).R.READY,
      saxigp5_awqos => s_axi_hp_in(3).AW.QOS, --[3:0]
      saxigp5_arqos => s_axi_hp_in(3).AR.QOS, --[3:0]

--resets using gpio
      pl_resetn0 => ps_out.FCLKRESET_N,
      --pl_resetn1 => open,
      --pl_resetn2 => open,
      --pl_resetn3 => open,

--For Clock buffering
--FCLK
      --pl_clk3 => ps_out.FCLK(3),
      --pl_clk2 => ps_out.FCLK(2),
      --pl_clk1 => ps_out.FCLK(1),
      pl_clk0 => ps_out.FCLK(0) --,
      );
end rtl;
