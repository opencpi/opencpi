../../../bias_param.rcc/target-1-linux-c6-x86_64/generics.vhd