-- THIS FILE WAS ORIGINALLY GENERATED ON Sat Apr  5 15:37:08 2014 EDT
-- BASED ON THE FILE: raw_test.xml
-- YOU *ARE* EXPECTED TO EDIT IT
-- This file initially contains the architecture skeleton for worker: raw_test

library IEEE; use IEEE.std_logic_1164.all; use ieee.numeric_std.all;
library ocpi; use ocpi.types.all; -- remove this to avoid all ocpi name collisions
architecture rtl of raw_test_worker is
begin
end rtl;
